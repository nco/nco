// Purpose: Generate a group file structure with common and non-common objects; pair of files are in_grp_1.cdl and in_grp_2.cdl
// Purpose: Pair of (different) files for 2 input file operators; pair of files are in_1.cdl and in_2.cdl
// Generate netCDF files with:
// ncgen -k netCDF-4 -b -o ~/nco/data/in_1.nc ~/nco/data/in_1.cdl
// ncgen -k netCDF-4 -b -o ~/nco/data/in_2.nc ~/nco/data/in_2.cdl

netcdf in_2 {
  dimensions:
  lon1=4;
  variables:
  float var1(lon1);
  data:
  var1=0,0,0,0;
} // end root group

