netcdf cf2 {
 // ncgen -k netCDF-4 -b -o ~/nco/data/cf2.nc ~/nco/data/cf2.cdl
 dimensions:
  lat=3;

 group: g1 {
  dimensions:
   lat=2;
  variables:
    float g1v1;
    g1v1:coordinates="/lat";
  data:
    g1v1=273.0;
  } // /g1

 group: g2 {
  dimensions:
    lat=2;
  variables:
    double lat(lat);
  data:
   lat=-90,90;
  } // /g2

} // end root group
