// Purpose: Generate test case for nces ensembles
// Generate netCDF files with:
// ncgen -k netCDF-4 -b -o ~/nco/data/in_grp_6.nc ~/nco/data/in_grp_6.cdl

netcdf in_grp_6 {

 group: cesm {

  group: cesm_01 {
  
   dimensions:
    lat=2;
    lon=4;
    time=unlimited; 
	
   variables:
    double time(time);
    float lat(lat);
    float lon(lon);
   
    float three_dmn_rec_var(time,lat,lon);
	
	data:
     lat=-90,90;
     lon=0,90,180,270;
     time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;

     three_dmn_rec_var=1, 2, 3, 4, 5, 6, 7, 8,
      9,10,11,12,13,14,15,16,
      17,18,19,20,21,22,23,24,
      25,26,27,28,29,30,31,32,
      33,34,35,36,37,38,39,40,
      41,42,43,44,45,46,47,48,
      49,50,51,52,53,54,55,56,
      57,58,59,60,61,62,63,64,
      65,66,67,68,69,70,71,72,
      73,74,75,76,77,78,79,80;
 
    } // cesm_01

  group: cesm_02 {
     
	
   dimensions:
    lat=2;
    lon=4;
    time=unlimited; 
	
   variables:
    double time(time);
    float lat(lat);
    float lon(lon);
   
    float three_dmn_rec_var(time,lat,lon);
	
	data:
     lat=-90,90;
     lon=0,90,180,270;
     time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;

     three_dmn_rec_var=1, 2, 3, 4, 5, 6, 7, 8,
      9,10,11,12,13,14,15,16,
      17,18,19,20,21,22,23,24,
      25,26,27,28,29,30,31,32,
      33,34,35,36,37,38,39,40,
      41,42,43,44,45,46,47,48,
      49,50,51,52,53,54,55,56,
      57,58,59,60,61,62,63,64,
      65,66,67,68,69,70,71,72,
      73,74,75,76,77,78,79,80;
 
    } // cesm_02
    
  } // cesm
  
} // root group
