// -*-C++-*-
// Purpose: CDL file to generate netCDF4 test file for vlen types

// Created: 20180413 based on buggy.cdl

// Usage:
// NB: ncgen arguments depend on version:
// "-k netCDF-4" for netCDF >= 3.6.3, "-k hdf5" for netCDF < 3.6.3
// "-k netCDF-4 classic model" for netCDF >= 3.6.3, "-k hdf5-nc3" for netCDF < 3.6.3
// ncgen -k netCDF-4 -b -o ~/nco/data/vlen.nc ~/nco/data/vlen.cdl
// scp ~/nco/data/vlen.cdl givre.ess.uci.edu:nco/data
// scp ~/nco/data/vlen.nc dust.ess.uci.edu:/var/www/html/nco
// scp dust.ess.uci.edu:/var/www/html/nco/vlen.nc ~/nco/data

netcdf vlen {

 types:
  // Declare all base-types of vlen's stored in file
  float(*) vlen_flt_t;
  int(*) vlen_int_t;
  short(*) vlen_sht_t;
  char(*) vlen_chr_t;
  uint64(*) vlen_uint64_t;
  string(*) vlen_sng_t; 
 dimensions:
  lat=2;
  lon=4;
  tm=10;  
  time=unlimited; 

 variables:
  int one;
  one:long_name="char attribute for one";

  float two;
  two:long_name="char attribute for two";
  
  vlen_flt_t vlen_flt_2D(lat,time);
  
  vlen_int_t vlen_int_scl;
  vlen_int_scl:long_name="vlen with base type integer";
  vlen_int_scl:number73=73;
  vlen_int_scl:_FillValue={-999}; // vlen data MUST BE enclosed in braces
  vlen_int_scl:number74=74;
  vlen_flt_t vlen_int_scl:vlen_att_flt_1D={1,2,3,4,5,6,7},{8,nanf,10};
  vlen_int_scl:flt_att_1D=1.0f,2.0f,3.0f,4.0f,5.0f,6.0f,7.0f,8.0f,nanf,10.0f;
  vlen_int_t vlen_int_scl:vlen_att_int_scl={1,2,3,4,5,6,7};
  vlen_int_t vlen_int_scl:vlen_att_int_1D={1,2,3,4,5,6,7},{8,9,10};
  vlen_sht_t vlen_int_scl:vlen_att_sht_1D={1,2,3,4,5,6,7},{8,9,10};
  vlen_int_scl:sht_att_1D=1s,2s,3s,4s,5s,6s,7s,8s,9s,10s;
  vlen_uint64_t vlen_int_scl:vlen_att_uint64_1D={1,2,3,4,5,6,7},{8,9,10};
  vlen_int_scl:uint64_att_1D=1ull,2ull,3ull,4ull,5ull,6ull,7ull,8ull,9ull,10ull;
  char vlen_int_scl:char_att="character attribute";
  float vlen_int_scl:flt_att=1.0;
  string vlen_int_scl:sng_att="string attribute";
  vlen_int_scl:_FillValue={-999};

  vlen_int_t vlen_int_1D(lat);
  vlen_int_1D:_FillValue={-999};

  vlen_int_t vlen_int_scl_mss_val_1D;
  vlen_int_scl_mss_val_1D:_FillValue={-999,-999}; // vlen data MUST BE enclosed in braces

  vlen_flt_t vlen_flt_scl;
  // 20180603: Investigate three _FillValue cases:
  // A. If _FillValue is not manually assigned, ncgen translates CDL underscores to default _FillValue of base type = 9.96921e+36 for floats, which is expected and seems correct 
  // B. If _FillValue is manually assigned, and CDL data section explicitly uses numeric value(s) (rather than an underscore) then ncgen correctly identifies that numeric values as the _FillValue.
  // C. For an underscore used in place of a single element within a VLEN, ncgen correctly uses default _FillValue of base type for the value of that element
  vlen_flt_scl:_FillValue={-999};

  vlen_flt_t vlen_flt_1D(lat);
  vlen_flt_1D:long_name="vlen with base type float";

  vlen_sng_t vlen_sng(lat);

  vlen_int_t three_dmn_var_vlen(tm,lat,lon);
  three_dmn_var_vlen:long_name="three dimensional record variable of type int";
  three_dmn_var_vlen:units="watt meter-2";
  three_dmn_var_vlen:_FillValue={-999};
  
 data:
  one=1;
  two=2;
  //  vlen_flt_scl={-999,17,18,19};
  // vlen_flt_scl={17,18,19};
  vlen_flt_scl=_;
  vlen_flt_2D={{1,2},{3,4}},{{5,6},{7,8}};
  vlen_flt_1D={17,18,19},{1,2,3,4,5,6,7,8,9,10};
  //vlen_int_scl={17,18,19};
  vlen_int_scl=_;
  vlen_int_1D=_,{1,2,3,4,5,6,7,8,9,10};
  vlen_int_scl_mss_val_1D=_;
  vlen_sng={"one","two","three"},{"four,five"};

  three_dmn_var_vlen= _, {2}, {3}, {4}, {5}, {6}, {7}, {8},
		     {9,9}, {10}, {11}, {12}, {13}, {14}, {15}, {16},
		     {17}, {18,18}, {19}, {20}, {21}, {22}, {23}, {24},
		     {25}, {26}, {27,27}, {28}, {29}, {30}, {31}, {32},
		     {33}, {34}, {35}, {36,36}, {37}, {38}, {39}, {40},
		     {41}, {42}, {43}, {44}, {45,45}, {46}, {47}, {48},
		     {49}, {50}, {51}, {52}, {53}, {54,54,54,54}, {55}, {56},
		     {57}, {58}, {59}, {60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75}, {61}, {62}, {63}, 
		     {65}, {66}, {67}, {68}, {69}, {70}, {71,62,73,74}, {72},
		     _, {74}, {75}, {76}, {77}, {78}, {79}, {80,81,82,83,84,85};

} // end root group
