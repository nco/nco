// -*-C++-*-
// Purpose: CDL file to generate netCDF4 test file for enum types

// Created: 20180413 based on buggy.cdl

// Usage:
// NB: ncgen arguments depend on version:
// "-k netCDF-4" for netCDF >= 3.6.3, "-k hdf5" for netCDF < 3.6.3
// "-k netCDF-4 classic model" for netCDF >= 3.6.3, "-k hdf5-nc3" for netCDF < 3.6.3
// ncgen -k netCDF-4 -b -o ~/nco/data/enum.nc ~/nco/data/enum.cdl
// scp ~/nco/data/enum.cdl givre.ess.uci.edu:nco/data
// scp ~/nco/data/enum.nc dust.ess.uci.edu:/var/www/html/nco
// scp dust.ess.uci.edu:/var/www/html/nco/enum.nc ~/nco/data

netcdf enum {

 // 20180413: types declarations must be first element in group, and appear before everything else. Where is this documented?
 types:
   ubyte enum enum_ubyte_t {Clear=0,Cumulonimbus=1,Stratus=2,Missing=128};
   short enum enum_sht_t {Small=-32000,Medium=0,Large=32767,missing_value=-32768};
   uint enum enum_uint_t {Greek_Καλημέρα=0,Japanese_キャク=1,Chinese_龥=3};
 // 20180522: Until today the base type of cargo was uint64. Changed it to uint because toolsUI 4.6.11 XML barfs on int64/uint64 enum because NcML lacks enum8 type. Once this changes can revert to uint64 (which works fine with C-library, NCO, and ncdump).
   uint64 enum cargo {bags\ of\ the\ best\ Sligo\ rags = 1000000, 
		      barrels\ of\ bones = 2000000, 
		      bails\ of\ old\ nanny\ goats\'\ tails = 3000000, 
		      barrels\ of\ stones = 4000000, dogs = 5000000, hogs = 6000000, 
		      barrels\ of\ porter = 7000000, 
		      sides\ of\ old\ blind\ horses\ hides = 8000000};
   int enum daysofWeekType { Monday = 1, Tuesday = 2, Wednesday = 3, Thursday= 4, Friday = 5, Saturday = 6, Sunday = 7 } ;

 dimensions:
   lat=2;
   lon=4;
   rec=8;

 variables:
   enum_ubyte_t cld_flg(lon);
   enum_ubyte_t cld_flg:_FillValue=Missing;

   enum_sht_t size(lon);
   enum_sht_t size:_FillValue=missing_value;

   enum_uint_t language(lon);
 
   cargo in_the_hold_of_the_Irish_Rover(lon);

   daysofWeekType days(lat, lon, rec);
 // 20180515: netCDF bug _FillValue must be a member otherwise default does not work see https://github.com/Unidata/netcdf-c/issues/982
   cargo in_the_hold_of_the_Irish_Rover:_FillValue=hogs;

 data:
   cld_flg=Stratus,_,Cumulonimbus,Clear;
   size=_,Small,Medium,Large;
   language=Chinese_龥,Japanese_キャク,Greek_Καλημέρα,Greek_Καλημέρα;
   in_the_hold_of_the_Irish_Rover=bags\ of\ the\ best\ Sligo\ rags,_,_,_;

 days= Monday, Tuesday,  Wednesday,  Thursday, Friday,  Saturday, Sunday, Monday,
       Monday, Tuesday,  Wednesday,  Thursday, Friday,  Saturday, Sunday, Monday,
       Monday, Tuesday,  Wednesday,  Thursday, Friday,  Saturday, Sunday, Monday,
       Monday, Tuesday,  Wednesday,  Thursday, Friday,  Saturday, Sunday, Monday,
       Monday, Tuesday,  Wednesday,  Thursday, Friday,  Saturday, Sunday, Monday,
       Monday, Tuesday,  Wednesday,  Thursday, Friday,  Saturday, Sunday, Monday,
       Monday, Tuesday,  Wednesday,  Thursday, Friday,  Saturday, Sunday, Monday,
       Monday, Tuesday,  Wednesday,  Thursday, Friday,  Saturday, Sunday, Monday,
       Monday, Tuesday,  Wednesday,  Thursday, Friday,  Saturday, Sunday, Monday,
       Monday, Tuesday,  Wednesday,  Thursday, Friday,  Saturday, Sunday, Monday;
 
} //end root group
