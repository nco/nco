// -*-C++-*-
// Purpose: File to test ncdismember
// Contains nested ensembles, metadata-only leaf groups, and "in-between data"
// Usage:
// ncgen -k netCDF-4 -b -o ~/nco/data/dsm.nc ~/nco/data/dsm.cdl
// ncdismember ~/nco/data/dsm.nc /data/zender/nco/tmp cf 1.5 > ~/foo.txt 2>&1

netcdf dsm {

  group: g1 {

  group: g1g1 {
      :metadata = "Leaf-group metadata";
    } // g1g1

  } // g1

  group: g2 {
    :metadata = "g2 group contains metadata and one variable but no shared dimensions";
  variables:
    float one;
    one:long_name="the loneliest number";
  data:
    one=1;
  } // g2

  group: g3 {
    :metadata = "g3 group contains metadata and one variable and one dimension";
  dimensions:
    lat=2;
  variables:
    float one_arr(lat);
    one_arr:long_name="the loneliest array";
  data:
    one_arr=1,1;
  } // g3

  group: g4 {
    :metadata = "g4 group contains one dimension, and one subgroup";
  dimensions:
    lat=2;
    group: g4g1 {
      :metadata = "g4g1 group contains one variable that depends on an inherited dimension";
    variables:
      float one_arr(lat);
      one_arr:long_name="the loneliest array";
    data:
      one_arr=1,1;
    } // g4g1

  } // g4

  group: g5 {
    :metadata = "g5 group contains one dimension, one variable (in-between) data and one subgroup";
  dimensions:
    lat=2;
  variables:
    float one_arr(lat);
    one_arr:long_name="the loneliest array";
    group: g5g1 {
      :metadata = "g5g1 group contains one variable that depends on an inherited dimension";
    variables:
      float one_arr(lat);
      one_arr:long_name="the loneliest array";
    data:
      one_arr=1,1;
    } // g5g1

  } // g5

  group: g6 {
    :metadata = "g6 group contains variables to test CF checkers";
  dimensions:
    time_like_2=2;
    time_like_3=2;
  variables:
    int period;
    period:units="second";
    period:long_name="length of time between successive orbits";
    byte time_like_1;
    time_like_1:units="ns";
    time_like_1:long_name="time";
    byte time_like_2(time_like_2);
    time_like_2:units="ns";
    time_like_2:long_name="time";
    byte time_like_3(time_like_3);
    time_like_3:calendar="none";
    time_like_3:units="ns";
    time_like_3:long_name="time";
    data:
    period=1;
    time_like_1=1b;
    time_like_2=1b,2b;
    time_like_3=1b,2b;
  } // g6

  group: cesm {

  group: cesm_01 {
      :Conventions = "CF-1.5";
      :history = "yada yada yada";
      :Scenario = "Historical";
      :Model = "CESM";
      :Realization = "1";

    dimensions:
      time=4;
    variables:
      float tas1(time);
      tas1:long_name="temperature";
      float tas2(time);
      tas2:long_name="temperature";
    data:
      tas1=272.1,272.1,272.1,272.1;
      tas2=272.1,272.1,272.1,272.1;
 
    } // cesm_01

  group: cesm_02 {
      :Conventions = "CF-1.5";
      :history = "yada yada yada";
      :Scenario = "Historical";
      :Model = "CESM";
      :Realization = "2";
      
    dimensions:
      time=4;
    variables:
      float tas1(time);
      tas1:long_name="temperature";
      float tas2(time);
      tas2:long_name="temperature";
    data:
      tas1=272.2,272.2,272.2,272.2;
      tas2=272.2,272.2,272.2,272.2;
      
    } // cesm_02
    
  } // cesm
  
 group: ecmwf {
    
  group: ecmwf_01 {
      :Conventions = "CF-1.5";
      :history = "yada yada yada";
      :Scenario = "Historical";
      :Model = "ECMWF";
      :Realization = "1";
      
    dimensions:
      time=4;
    variables:
      float tas1(time);
      tas1:long_name="temperature";
      float tas2(time);
      tas2:long_name="temperature";
    data:
      tas1=273.1,273.1,273.1,273.1;
      tas2=273.1,273.1,273.1,273.1;
      
    } // ecmwf_01
    
  group: ecmwf_02 {
      :Conventions = "CF-1.5";
      :history = "yada yada yada";
      :Scenario = "Historical";
      :Model = "ECMWF";
      :Realization = "2";
      
    dimensions:
      time=4;
    variables:
      float tas1(time);
      tas1:long_name="temperature";
      float tas2(time);
      tas2:long_name="temperature";      
    data:
      tas1=273.2,273.2,273.2,273.2;
      tas2=273.2,273.2,273.2,273.2;
    } // ecmwf_02

  } // ecmwf

} // root group
