// $Header: /data/zender/nco_20150216/nco/bm/gne_exp.cdl,v 1.3 2005-04-19 21:19:49 mangalam Exp $
// Purpose: CDL file to generate a netCDF file that approximates a gene expression data set.

// Usage:
// Create ge.nc from ge.cdl on a beefy 64-bit computer
// ncgen -b -o ge.nc ge.cdl

// On small-RAM machines, create 50MB file with multiple simple variables
// ncap -D 3 -O -s "wvl_1e8[wvl_1e8]=1.0f" ~/nco/data/big.nc ${DATA}/tmp/big.nc

// Valid CDF/netCDF files need not have any defined variable or data

// Use ncap LHS-casting to define variables with big dimensions
netcdf mlw_gene_ex{
dimensions:
//replicates per cell
    rep=3;
//treatment per cell
    treat=2;
//number of cell types tested
    cell=4;
//# of parameters per 'gene' or ge_atom)
    params=10;
//# of genes thingies tested for - let it grow
    ge_atoms=unlimited;
    
variables:
    double ge_atoms(ge_atoms);
    double rep(rep);
    double treat(treat);
    double cell(cell);
    double params(params);
    float base(ge_atoms,rep,treat,cell,params);
data:
}
