// -*-C++-*-
// Purpose: 
// ncpdq tests
// Generate netCDF files with:
// ncgen -k netCDF-4  -b -o ~/nco/data/in_grp_8.nc ~/nco/data/in_grp_8.cdl

netcdf in_grp_8 {
 group: g1 { 
   dimensions:
    lat=2;
    lon=3;
    time=unlimited;
    variables:
    float lat(lat);
    float lon(lon);
    double time(time);
    float snd(time,lat,lon);
    data:
    lat=0,1;
    lon=0,1,2;
    time=0,1;
    snd=0,1,2,3,4,5,6,7,8,9,10,11;
  } // end g1
  
  group: g2 { 
   dimensions:
    lat=2;
    lon=3;
    time=unlimited;
    variables:
    float lat(lat);
    float lon(lon);
    double time(time);
    float snd(time,lat,lon);
    data:
    lat=0,1;
    lon=0,1,2;
    time=0,1;
    snd=0,1,2,3,4,5,6,7,8,9,10,11;
  } // end g2
 
} // root group
