// ncgen -b -o ~/nco/data/nco_gsl.nc ~/nco/data/nco_gsl.cdl

netcdf nco_gsl {
//purpose: test nco_gsl_fit_linear()
//usage: ncap2 -O -S ~/nco/data/nco_gsl.nco ~/nco/data/nco_gsl.nc out.nc      
//case 1; vx,vy   double arrays with no fill value and dim=N
//case 2; fx,fy   double arrays one fill value in fy and dim=N
//case 3; vxr,vyr double arrays with no fill value and dim=N-1, index a fill value case 2 removed
//case 2 and case 3 must return the same values for: &c0,&c1,&cov00,&cov01,&cov11,&sumsq
	dimensions:
	dim=4;
	dimr=3;
	variables:
	double vx(dim);
	double vy(dim);
	double fx(dim);
	double fy(dim);
	fy:_FillValue = -99.0;
	double vxr(dimr);
	double vyr(dimr);
	data:
	vx=2.0,3.0,2.0,3.0;
	vy=4.0,6.0,6.0,8.0;
	fx=2.0,3.0,2.0,3.0;
	fy=4.0,-99.0,6.0,8.0;
	vxr=2.0,2.0,3.0;
	vyr=4.0,6.0,8.0;
}
