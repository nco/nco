// ncgen -k netCDF-4 -b -o ~/nco/data/cmip5.nc ~/nco/data/cmip5.cdl

netcdf cmip5 {
  :Conventions = "CF-2.x";
  :history = "yada yada yada";
  :Scenario = "RCP 8.5";

  group: cesm { 
  dimensions:
  time=unlimited;
  variables:
  float tas(time);
  :Model = "CESM";
  data:
  tas=272,272,272,272;
  } // end cesm
  
  group: ecmwf { 
  dimensions:
  time=unlimited;
  variables:
  float tas(time);
  :Model = "ECMWF";
  data:
  tas=273,273,273,273;
  } // end ecmwf
  
  group: giss { 
  dimensions:
  time=unlimited;
  variables:
  float tas(time);
  :Model = "GISS";
  data:
  tas=274,274,274,274;
  } // end gfdl

} // end root group
