netcdf split {
dimensions:
	time = UNLIMITED ; // (36 currently)
	ncol = 101 ;
	nbnd = 2 ;
variables:
	float AODVIS(time, ncol) ;
		AODVIS:_FillValue = 1.e+36f ;
		AODVIS:missing_value = 1.e+36f ;
		AODVIS:units = "" ;
		AODVIS:long_name = "Aerosol optical depth 550 nm" ;
		AODVIS:cell_methods = "time: mean" ;
	double area(ncol) ;
	double lat(ncol) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
	double lon(ncol) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nbnd) ;
		time_bnds:long_name = "time interval endpoints" ;

// global attributes:
		:np = 4 ;
		:ne = 30 ;
		:Conventions = "CF-1.0" ;
		:source = "CAM" ;
		:case = "famipc5_ne30_v0.3_00003" ;
		:title = "UNSET" ;
		:logname = "mbranst" ;
		:host = "nid02435" ;
		:Version = "$Name$" ;
		:revision_Id = "$Id$" ;
		:initial_file = "/scratch2/scratchdirs/mbranst/acme_scratch/inputdata/ne30_gx1.F1850c5d.cam.i.0006-01-01-00000.nc" ;
		:topography_file = "/project/projectdirs/ccsm1/inputdata/atm/cam/topo/USGS-gtopo30_ne30np4_16xdel2-PFC-consistentSGH.nc" ;
		:NCO = "\"4.6.0\"" ;
		:nco_openmp_thread_number = 1 ;
data:

 AODVIS =
  0.1954915, 0.2052418, 0.2055524, 0.1982304, 0.2047635, 0.2120854, 0.184495, 
    0.193814, 0.1982379, 0.1796773, 0.1873291, 0.1900486, 0.2092419, 
    0.2124223, 0.2095956, 0.2165151, 0.2197439, 0.2198535, 0.2026321, 
    0.210454, 0.2129825, 0.1927225, 0.1985276, 0.1994585, 0.2075444, 
    0.2046486, 0.2036938, 0.2174332, 0.2119768, 0.2074966, 0.2119771, 
    0.2063783, 0.2007158, 0.1984009, 0.1980032, 0.1993936, 0.2027589, 
    0.1959963, 0.1937612, 0.2026193, 0.1953114, 0.1911157, 0.1940382, 
    0.1907044, 0.1884757, 0.2003334, 0.1979246, 0.1983925, 0.1914183, 
    0.1890862, 0.1885663, 0.1891981, 0.1897797, 0.1897665, 0.1884398, 
    0.1926364, 0.1953603, 0.2011434, 0.2019434, 0.2036232, 0.1881192, 
    0.1881149, 0.1857819, 0.1922142, 0.1915971, 0.1921426, 0.1979958, 
    0.198307, 0.196068, 0.2012686, 0.2007759, 0.2006028, 0.1859224, 
    0.1863353, 0.1868506, 0.1925839, 0.1933768, 0.1940954, 0.1969706, 
    0.1940695, 0.1951418, 0.199446, 0.196628, 0.1943224, 0.188907, 0.1917336, 
    0.1935624, 0.195038, 0.1972754, 0.1976926, 0.1923693, 0.1948078, 
    0.1949104, 0.1940187, 0.194156, 0.1961968, 0.1962795, 0.1968865, 
    0.1959289, 0.200077, 0.1979352,
  0.08774699, 0.08743263, 0.08813152, 0.08697822, 0.08712716, 0.08697484, 
    0.08066922, 0.08181216, 0.08227495, 0.07723534, 0.08017638, 0.08140094, 
    0.09060917, 0.09402835, 0.09687552, 0.08742309, 0.0918293, 0.09480345, 
    0.08381522, 0.08884465, 0.09221447, 0.0819945, 0.08621505, 0.09087382, 
    0.09871756, 0.1039915, 0.1066364, 0.09834164, 0.1046, 0.1087259, 
    0.09643233, 0.1029484, 0.1073058, 0.09439981, 0.1007063, 0.1042427, 
    0.1086272, 0.1132357, 0.1164022, 0.1122138, 0.1168153, 0.1192327, 
    0.1101353, 0.1146111, 0.1164792, 0.10632, 0.1101103, 0.1108131, 
    0.1174577, 0.1194424, 0.1198301, 0.1208031, 0.1236182, 0.1253759, 
    0.1161827, 0.1195217, 0.121555, 0.1105978, 0.1127567, 0.1138001, 
    0.1241897, 0.129181, 0.1299398, 0.1274792, 0.1320326, 0.1333827, 
    0.1222774, 0.1241962, 0.1269779, 0.1142067, 0.1131517, 0.1144032, 
    0.1315697, 0.1317602, 0.132011, 0.1356063, 0.1343876, 0.1365362, 
    0.1273904, 0.1286372, 0.1312875, 0.1174474, 0.1185959, 0.1207921, 
    0.1325194, 0.1315188, 0.1314559, 0.1350825, 0.1362105, 0.1351408, 
    0.1304566, 0.1318385, 0.1342105, 0.1245243, 0.1285835, 0.1316005, 
    0.1317033, 0.1362245, 0.1395495, 0.1373214, 0.1429455,
  0.1739239, 0.1729402, 0.1719707, 0.1711836, 0.174391, 0.1745256, 0.1603207, 
    0.157661, 0.1594325, 0.1611351, 0.1577098, 0.1590508, 0.1724134, 
    0.1728314, 0.1737903, 0.1757511, 0.176421, 0.1767885, 0.1627198, 
    0.170582, 0.1744228, 0.164528, 0.1702799, 0.1709895, 0.1761124, 
    0.1808682, 0.1801839, 0.1775861, 0.177875, 0.1742473, 0.1755064, 
    0.165073, 0.1578238, 0.1693932, 0.1585429, 0.1538348, 0.1803929, 
    0.1798392, 0.1750582, 0.1709813, 0.1658825, 0.1617512, 0.1529435, 
    0.148134, 0.14108, 0.1465365, 0.1392745, 0.1349678, 0.1716387, 0.1645602, 
    0.1612926, 0.1581703, 0.1528563, 0.1519293, 0.1396111, 0.1401398, 
    0.1405889, 0.1335033, 0.1348822, 0.1368755, 0.1606339, 0.1534593, 
    0.1538814, 0.1529485, 0.152769, 0.1529377, 0.1432214, 0.1452122, 
    0.1481796, 0.1389131, 0.137797, 0.1354714, 0.15597, 0.1617808, 0.1656674, 
    0.1564982, 0.1605673, 0.1622002, 0.1489572, 0.1474354, 0.1448696, 
    0.1318119, 0.1297729, 0.1316136, 0.1686257, 0.1727131, 0.1759136, 
    0.1636261, 0.165663, 0.1689182, 0.1458476, 0.1497804, 0.1498627, 
    0.1353435, 0.1402377, 0.1444481, 0.1779456, 0.1853191, 0.1852839, 
    0.1681498, 0.1714406,
  0.1786167, 0.1873076, 0.194791, 0.1864717, 0.1993225, 0.206763, 0.1901386, 
    0.1990162, 0.2026069, 0.1908278, 0.193333, 0.1941527, 0.2006553, 0.2057, 
    0.2014703, 0.2170719, 0.2169071, 0.2115936, 0.2038641, 0.2006001, 
    0.1951292, 0.1940284, 0.1871726, 0.1834531, 0.198143, 0.1883013, 
    0.1789255, 0.203945, 0.194141, 0.1842929, 0.1911463, 0.1842547, 0.179635, 
    0.1815618, 0.179608, 0.1766685, 0.1752679, 0.1709059, 0.1707577, 
    0.1767845, 0.1709922, 0.1708429, 0.1759156, 0.1752726, 0.1783778, 
    0.1749188, 0.177655, 0.1779721, 0.1725561, 0.174211, 0.174641, 0.1754592, 
    0.1814622, 0.1812453, 0.1798575, 0.1822189, 0.177544, 0.1792191, 
    0.1805906, 0.1779069, 0.1763419, 0.1754508, 0.1706967, 0.1789466, 
    0.1694007, 0.1647493, 0.1712515, 0.1614626, 0.1580704, 0.1743896, 
    0.1646255, 0.1600677, 0.1648719, 0.1568906, 0.1547807, 0.1599964, 
    0.1554217, 0.1554395, 0.1565195, 0.1581038, 0.1590432, 0.162646, 
    0.1611406, 0.1604452, 0.1528743, 0.1513192, 0.1497111, 0.1586315, 
    0.1562136, 0.1562016, 0.1655106, 0.1636323, 0.1619447, 0.160639, 
    0.1601082, 0.1592852, 0.1492148, 0.1500751, 0.1525081, 0.1563363, 0.160644,
  0.1510869, 0.1542146, 0.156989, 0.1632795, 0.1673208, 0.1679074, 0.1927984, 
    0.2025148, 0.203211, 0.2143254, 0.21573, 0.2130025, 0.1603853, 0.1657471, 
    0.1676381, 0.1704904, 0.1730234, 0.1732247, 0.2015578, 0.1927796, 
    0.1877322, 0.208733, 0.2018969, 0.1967425, 0.1700829, 0.1717525, 
    0.1729111, 0.1740752, 0.1770962, 0.1760429, 0.1853302, 0.1847549, 
    0.1870149, 0.1945629, 0.1952988, 0.1985721, 0.1748789, 0.1819272, 
    0.1849024, 0.1767615, 0.1795637, 0.1793738, 0.1887766, 0.1918996, 
    0.1945476, 0.1997209, 0.2044196, 0.2060402, 0.188743, 0.1842763, 
    0.1748654, 0.1774349, 0.1770387, 0.1749263, 0.1968132, 0.199715, 
    0.1992591, 0.2058188, 0.2077636, 0.2106776, 0.170015, 0.1579867, 
    0.153783, 0.1710836, 0.1675183, 0.1664319, 0.1997712, 0.1993994, 
    0.1991671, 0.2138371, 0.2140347, 0.2106524, 0.1581412, 0.1591951, 
    0.1613065, 0.1704873, 0.1677732, 0.166469, 0.1961351, 0.1909115, 
    0.1870097, 0.2027994, 0.1919652, 0.1877802, 0.1588414, 0.1552486, 
    0.1553995, 0.1674631, 0.1674751, 0.168565, 0.1866269, 0.1858682, 
    0.1832919, 0.1861531, 0.187217, 0.1871001, 0.1577048, 0.165372, 
    0.1682718, 0.16802, 0.1742394,
  0.1906363, 0.1901704, 0.1875623, 0.2025749, 0.206433, 0.2005123, 0.2170124, 
    0.2204212, 0.2193098, 0.2362882, 0.2321109, 0.2297994, 0.1846904, 
    0.181544, 0.1781296, 0.19502, 0.1966698, 0.1865541, 0.2076659, 0.2046331, 
    0.2122996, 0.2244332, 0.2236025, 0.2221671, 0.1726549, 0.1683958, 
    0.1630023, 0.1866049, 0.1762094, 0.1740675, 0.2065514, 0.2078829, 
    0.2042466, 0.2239724, 0.2190723, 0.2153239, 0.1609292, 0.1569534, 
    0.1546557, 0.1699765, 0.1666802, 0.1687745, 0.2048534, 0.1955038, 
    0.1923232, 0.2117693, 0.2075251, 0.2058202, 0.1509489, 0.1497327, 
    0.1481774, 0.1681512, 0.1666452, 0.1628895, 0.1905132, 0.1884256, 
    0.1891769, 0.2044083, 0.2005369, 0.2022443, 0.1481222, 0.1447443, 
    0.1471749, 0.1592498, 0.1619628, 0.1635137, 0.1870604, 0.1917661, 
    0.192659, 0.2035804, 0.2065762, 0.2076468, 0.1453881, 0.1448493, 
    0.1440915, 0.1644577, 0.165576, 0.1662327, 0.1950034, 0.1953014, 
    0.1949191, 0.207452, 0.2062996, 0.2137531, 0.146671, 0.1498499, 
    0.1521496, 0.1694918, 0.1763436, 0.1811759, 0.2067915, 0.2116499, 
    0.2167345, 0.2138439, 0.2262517, 0.2315412, 0.1571211, 0.1640163, 
    0.1674957, 0.1874029, 0.1945786,
  0.1896786, 0.1918914, 0.1892491, 0.1962431, 0.2014005, 0.1992956, 
    0.2048586, 0.2066852, 0.2034762, 0.2082825, 0.2001792, 0.1949693, 
    0.1885221, 0.1902647, 0.1890659, 0.1961279, 0.1928118, 0.1887126, 
    0.199409, 0.1938328, 0.1902045, 0.1916712, 0.1888143, 0.1893841, 
    0.190686, 0.1909313, 0.1862512, 0.1912346, 0.1930633, 0.1907808, 
    0.1902959, 0.1921044, 0.1961961, 0.1935471, 0.1970171, 0.1975437, 
    0.1806876, 0.1817406, 0.1835687, 0.1862947, 0.1878512, 0.190567, 
    0.1982914, 0.1967019, 0.1975832, 0.2016835, 0.199562, 0.1941278, 
    0.1900091, 0.1964789, 0.1986384, 0.1920092, 0.1933239, 0.1931775, 
    0.1966315, 0.1903583, 0.183803, 0.1900206, 0.1853285, 0.1880271, 
    0.1987904, 0.1971742, 0.1927225, 0.1930726, 0.1922454, 0.1947364, 
    0.184542, 0.1896671, 0.1896102, 0.1912159, 0.1969684, 0.1913841, 
    0.1929263, 0.1847612, 0.1800319, 0.1909867, 0.1811586, 0.1714433, 
    0.1848235, 0.1768371, 0.173429, 0.1873626, 0.1790878, 0.1723381, 
    0.1759883, 0.168194, 0.1602721, 0.1666408, 0.1649366, 0.1626477, 
    0.1664855, 0.1602642, 0.1621723, 0.168886, 0.1638036, 0.1644865, 
    0.1601189, 0.1610846, 0.1612729, 0.1605711, 0.162232,
  0.2119588, 0.2176632, 0.2208682, 0.2152513, 0.2200734, 0.2240904, 
    0.2090581, 0.2107005, 0.2110124, 0.1987567, 0.2040146, 0.2046128, 
    0.2212195, 0.2174118, 0.2079995, 0.2229085, 0.2193937, 0.2159309, 
    0.2093493, 0.2101333, 0.2076997, 0.2052733, 0.2060551, 0.2072342, 
    0.2007361, 0.1909193, 0.1855097, 0.2077152, 0.1959265, 0.1881483, 
    0.20602, 0.2013719, 0.2005085, 0.2065096, 0.204934, 0.205859, 0.1844421, 
    0.1793746, 0.1768478, 0.1857276, 0.1854429, 0.1833152, 0.201065, 
    0.2031028, 0.2054031, 0.207064, 0.2125163, 0.2071044, 0.1746369, 
    0.1744489, 0.1762774, 0.1819557, 0.1840626, 0.185436, 0.2030785, 
    0.1988732, 0.1957376, 0.2078757, 0.2054155, 0.2026137, 0.1730461, 
    0.1723439, 0.1704763, 0.1824181, 0.1783503, 0.1802525, 0.1946535, 
    0.190704, 0.1911389, 0.2049982, 0.2037122, 0.2029213, 0.1697549, 
    0.1707603, 0.1701994, 0.1782067, 0.1799704, 0.1797967, 0.1904994, 
    0.18754, 0.1863115, 0.2003481, 0.1938203, 0.1926307, 0.1702934, 
    0.1698078, 0.1666698, 0.1795557, 0.178874, 0.1780438, 0.1881538, 
    0.1861796, 0.1829003, 0.1912631, 0.1895325, 0.1878059, 0.1681777, 
    0.1660794, 0.167106, 0.1789467, 0.1760756,
  0.1286334, 0.1269895, 0.127767, 0.1361609, 0.1354878, 0.1336268, 0.1465011, 
    0.1461069, 0.1402656, 0.1523714, 0.140247, 0.1372345, 0.1294348, 
    0.1283572, 0.1273577, 0.1334204, 0.1337974, 0.1340785, 0.1346631, 
    0.1310677, 0.1303914, 0.1363534, 0.1345273, 0.1342929, 0.1284832, 
    0.130027, 0.1312707, 0.1321506, 0.1340037, 0.1374296, 0.1303741, 
    0.1337655, 0.1365032, 0.1337021, 0.1340505, 0.1360545, 0.1344812, 
    0.1397676, 0.1411705, 0.1385749, 0.1422145, 0.1454634, 0.1372489, 
    0.1379296, 0.1394332, 0.1368502, 0.1394547, 0.1405112, 0.142928, 
    0.145283, 0.1440065, 0.1517887, 0.1514257, 0.1480746, 0.1405668, 
    0.1414474, 0.1392117, 0.14344, 0.1455315, 0.143189, 0.1420373, 0.1403603, 
    0.1400274, 0.1428212, 0.1386795, 0.1377767, 0.1389547, 0.1367873, 
    0.1389611, 0.1434318, 0.1434912, 0.1433651, 0.1392526, 0.1372387, 
    0.1316812, 0.1398527, 0.1362854, 0.1324909, 0.140595, 0.141123, 
    0.1401738, 0.1436628, 0.1457977, 0.1444397, 0.1294797, 0.1272952, 
    0.1283476, 0.1290243, 0.132112, 0.1339472, 0.1403411, 0.1439678, 
    0.1451737, 0.1451481, 0.1477971, 0.1471629, 0.1284245, 0.1340864, 
    0.1365195, 0.1384986, 0.1421767,
  0.1299628, 0.1294229, 0.1274931, 0.1345598, 0.1340972, 0.1325774, 
    0.1379275, 0.141089, 0.1393437, 0.1387298, 0.1412361, 0.1417763, 
    0.1283337, 0.1257687, 0.1237329, 0.1303241, 0.1293273, 0.1273175, 
    0.1368629, 0.1368748, 0.137399, 0.1407822, 0.1449397, 0.1426928, 
    0.1224963, 0.1217772, 0.1230937, 0.1249061, 0.1243884, 0.127071, 
    0.1357506, 0.1302515, 0.1255872, 0.1391151, 0.1289692, 0.1258496, 
    0.1265729, 0.1261442, 0.1295586, 0.1275589, 0.128249, 0.1298158, 
    0.1227465, 0.1242012, 0.1295258, 0.1239649, 0.1292922, 0.1390608, 
    0.1301167, 0.1319485, 0.1314989, 0.1323018, 0.135418, 0.1360931, 0.13685, 
    0.148744, 0.151734, 0.1489494, 0.1559564, 0.1586595, 0.1302561, 
    0.1306875, 0.1316861, 0.1348991, 0.1367945, 0.137563, 0.1534979, 
    0.1527037, 0.1522826, 0.159484, 0.1605415, 0.1575736, 0.1286758, 
    0.1246191, 0.1229084, 0.135054, 0.1334736, 0.1347913, 0.1497687, 
    0.1463766, 0.1484456, 0.1524964, 0.147383, 0.1415917, 0.1253459, 
    0.1306985, 0.1343014, 0.1380304, 0.1402359, 0.1408973, 0.1472926, 
    0.142153, 0.1399773, 0.138021, 0.1320983, 0.1306829, 0.1366407, 
    0.1398129, 0.1399482, 0.1436093, 0.141966,
  0.146344, 0.142248, 0.1393117, 0.1552604, 0.1531578, 0.1497421, 0.1563542, 
    0.158169, 0.1598406, 0.1535019, 0.1556785, 0.1577791, 0.1405883, 
    0.1488269, 0.1508076, 0.1517251, 0.1560772, 0.1619961, 0.1598524, 
    0.1668183, 0.1677451, 0.1593428, 0.164622, 0.1669476, 0.1523084, 0.15468, 
    0.1526962, 0.1635156, 0.1668611, 0.1685837, 0.1705939, 0.1744903, 
    0.1756771, 0.1644497, 0.1675043, 0.1689485, 0.1493731, 0.1463022, 
    0.1438671, 0.1696408, 0.1631103, 0.1638779, 0.1800926, 0.1868232, 
    0.1833488, 0.1742091, 0.1793512, 0.1798557, 0.1422958, 0.1377194, 
    0.1345088, 0.1606339, 0.1543148, 0.1494279, 0.1831117, 0.1813686, 
    0.1768945, 0.1813985, 0.1805276, 0.1794018, 0.1292731, 0.1276147, 
    0.126546, 0.1450379, 0.1438734, 0.1430462, 0.1741115, 0.1730857, 
    0.1764767, 0.1782845, 0.1786447, 0.1749635, 0.1269091, 0.1283551, 
    0.1301016, 0.1424581, 0.1450208, 0.1427712, 0.171021, 0.1654073, 
    0.1641171, 0.1747841, 0.1729056, 0.1682506, 0.1317082, 0.1303201, 
    0.1263227, 0.1443875, 0.1403969, 0.1363788, 0.1624428, 0.1551939, 
    0.1524396, 0.1650937, 0.1575785, 0.1571647, 0.1248747, 0.123309, 
    0.1232975, 0.1350061, 0.1329321,
  0.1755102, 0.1782824, 0.1814537, 0.1732881, 0.1765223, 0.1797348, 
    0.1697965, 0.1716152, 0.1735759, 0.1708749, 0.172013, 0.1716569, 
    0.184084, 0.1849064, 0.1850084, 0.1815074, 0.1810918, 0.1784322, 
    0.1749404, 0.1728542, 0.1660836, 0.1695973, 0.1634995, 0.1627289, 
    0.182243, 0.1759662, 0.1747504, 0.1755952, 0.1722731, 0.1706973, 
    0.1660955, 0.1647148, 0.1645323, 0.1583723, 0.1584442, 0.1574573, 
    0.1738243, 0.1744748, 0.1735976, 0.170867, 0.1720889, 0.1713889, 
    0.1650033, 0.1641487, 0.1615691, 0.1557691, 0.1532708, 0.1506609, 
    0.1730418, 0.1679271, 0.1627403, 0.1694104, 0.1623394, 0.156324, 
    0.1572356, 0.1524252, 0.1497952, 0.1495337, 0.14782, 0.1475905, 
    0.1577343, 0.1518547, 0.1485603, 0.151631, 0.1481112, 0.1495731, 
    0.1486705, 0.1479519, 0.1477144, 0.1469421, 0.1447637, 0.1441316, 
    0.148768, 0.1506405, 0.1511921, 0.1493118, 0.1517575, 0.1535962, 
    0.1478382, 0.146755, 0.1478933, 0.1433997, 0.1424003, 0.1417823, 
    0.1537059, 0.156788, 0.1595886, 0.1553896, 0.1575987, 0.1592122, 0.14973, 
    0.1535225, 0.1557317, 0.1481648, 0.1546776, 0.1572393, 0.1608133, 
    0.1618119, 0.1613342, 0.1591998, 0.1599037,
  0.139913, 0.1412289, 0.1455513, 0.1396898, 0.1435158, 0.1453746, 0.1463682, 
    0.1543897, 0.1567084, 0.1488611, 0.1526124, 0.1515827, 0.1498866, 
    0.1587924, 0.1638683, 0.1478017, 0.1554752, 0.1599506, 0.1573369, 
    0.158221, 0.1601354, 0.1523053, 0.1529154, 0.1535422, 0.1658488, 
    0.1716795, 0.1688759, 0.1647966, 0.1708144, 0.1736228, 0.1628351, 
    0.1701769, 0.1740719, 0.1555968, 0.1605071, 0.1639858, 0.165073, 
    0.1609458, 0.1570887, 0.1733034, 0.1754312, 0.174106, 0.1761086, 
    0.180278, 0.1807026, 0.1690371, 0.1715597, 0.1735135, 0.1529972, 
    0.1491329, 0.1452413, 0.1704442, 0.1661207, 0.1627326, 0.1784918, 
    0.1776706, 0.1736342, 0.173457, 0.1697119, 0.1692021, 0.1438615, 
    0.1433771, 0.1408377, 0.1599263, 0.1545115, 0.1549845, 0.1704183, 
    0.1652213, 0.1649592, 0.1668992, 0.1686076, 0.1720167, 0.1408773, 
    0.143125, 0.1423426, 0.1523266, 0.1515496, 0.152986, 0.1650627, 
    0.1655363, 0.1645259, 0.171628, 0.1737596, 0.1745078, 0.1426373, 
    0.1454382, 0.1491868, 0.1541699, 0.1574278, 0.1583546, 0.168814, 
    0.1652257, 0.1593018, 0.1736458, 0.1679257, 0.1633575, 0.1511276, 
    0.1509706, 0.1503545, 0.1592737, 0.1570367,
  0.1246863, 0.1219536, 0.1190693, 0.1254627, 0.1242086, 0.1250418, 
    0.1255953, 0.1275962, 0.1277172, 0.125637, 0.1281339, 0.1270378, 
    0.1196316, 0.1160785, 0.1148444, 0.1260579, 0.1257013, 0.1256686, 
    0.1269731, 0.1279412, 0.1275063, 0.1273239, 0.1279111, 0.1283612, 
    0.1137424, 0.1128109, 0.1135152, 0.1258531, 0.124796, 0.1229969, 
    0.1284424, 0.1306434, 0.1328965, 0.1276713, 0.1271854, 0.127332, 
    0.1134498, 0.1130523, 0.1143744, 0.1231111, 0.1248598, 0.1247131, 
    0.1345185, 0.1356363, 0.1344033, 0.129937, 0.130238, 0.1296404, 
    0.1142002, 0.1173661, 0.1196253, 0.1246305, 0.1247103, 0.12595, 0.133165, 
    0.1293872, 0.1263612, 0.1306048, 0.1269332, 0.1248906, 0.1234029, 
    0.1297777, 0.1319967, 0.1270217, 0.1287481, 0.1298174, 0.1254088, 
    0.1243806, 0.1233314, 0.1230178, 0.124957, 0.1239709, 0.1349693, 
    0.1414731, 0.1424994, 0.1305704, 0.1315547, 0.1321315, 0.1223826, 
    0.1238686, 0.1242745, 0.1270712, 0.1288312, 0.1327871, 0.1432531, 
    0.1444277, 0.1453653, 0.1316171, 0.1340172, 0.1343308, 0.1268829, 
    0.1317597, 0.1342965, 0.1356966, 0.1389286, 0.1411946, 0.1464154, 
    0.1480325, 0.1483928, 0.1361819, 0.1413696,
  0.160341, 0.1635033, 0.1621206, 0.1515452, 0.1585005, 0.1614555, 0.1398125, 
    0.1423866, 0.1456765, 0.1396807, 0.139869, 0.140501, 0.1608388, 
    0.1609773, 0.1592907, 0.1621868, 0.1657887, 0.1668044, 0.1475483, 
    0.1514947, 0.1539889, 0.1411643, 0.1427867, 0.1441789, 0.1590194, 
    0.1573306, 0.1560811, 0.1664279, 0.1654406, 0.161945, 0.155193, 
    0.1538208, 0.1558266, 0.1454617, 0.1457111, 0.1464898, 0.1561266, 
    0.1546205, 0.1530069, 0.1604971, 0.1599716, 0.1587257, 0.1572253, 
    0.1547799, 0.1563955, 0.1479519, 0.1481985, 0.1510885, 0.1519727, 
    0.153555, 0.153074, 0.1562887, 0.1563622, 0.1575526, 0.1564805, 
    0.1550865, 0.1581646, 0.150941, 0.1534169, 0.1538319, 0.1540512, 
    0.1600211, 0.1630145, 0.1586583, 0.159132, 0.1585571, 0.159025, 
    0.1616082, 0.1572852, 0.1535651, 0.1535514, 0.1523865, 0.16494, 
    0.1675206, 0.162421, 0.1588283, 0.1540163, 0.150922, 0.1515824, 
    0.1472509, 0.1467513, 0.1512851, 0.1503641, 0.1486479, 0.1594772, 
    0.1596295, 0.1619115, 0.1486044, 0.1501469, 0.1547556, 0.1452666, 
    0.1414726, 0.1406678, 0.1460992, 0.139055, 0.1331514, 0.1642474, 
    0.1722728, 0.1703433, 0.157058, 0.158688,
  0.2219688, 0.2192966, 0.218588, 0.2278748, 0.2287727, 0.2268884, 0.2317646, 
    0.242741, 0.2434133, 0.2411369, 0.2510195, 0.2544318, 0.213603, 
    0.2101426, 0.2105355, 0.2253622, 0.223389, 0.2198058, 0.2472358, 
    0.2482178, 0.2502292, 0.2557815, 0.2563511, 0.2557927, 0.2095963, 
    0.2095486, 0.2101364, 0.2169804, 0.213447, 0.2082549, 0.251557, 
    0.2455387, 0.2386892, 0.2533324, 0.2465655, 0.2405316, 0.2056717, 
    0.1949571, 0.1913736, 0.207105, 0.2046446, 0.2040785, 0.2327742, 
    0.2237252, 0.2179521, 0.233891, 0.2224127, 0.2150826, 0.1896309, 
    0.1904342, 0.1875363, 0.205963, 0.2023262, 0.2032399, 0.2127466, 
    0.2095153, 0.2096834, 0.2132701, 0.2085732, 0.2064312, 0.185988, 
    0.1858601, 0.1831141, 0.2041567, 0.2011562, 0.1985588, 0.2100198, 
    0.2120034, 0.2087582, 0.208389, 0.2103929, 0.2097145, 0.1810902, 
    0.1777561, 0.1766852, 0.1945111, 0.1896358, 0.1884039, 0.2032826, 
    0.1960589, 0.196144, 0.2109251, 0.2105203, 0.2097526, 0.1750808, 
    0.1778845, 0.1771683, 0.1862403, 0.1858459, 0.1862284, 0.194868, 
    0.1928691, 0.1948864, 0.2109767, 0.2136056, 0.2148038, 0.1746529, 
    0.1728472, 0.1708699, 0.1868666, 0.185789,
  0.2351467, 0.2232926, 0.2187398, 0.2140746, 0.2072348, 0.2054752, 
    0.1987498, 0.1946953, 0.1908217, 0.206033, 0.2007624, 0.1971389, 
    0.2156579, 0.2155334, 0.2131321, 0.2041002, 0.207699, 0.2126335, 
    0.1915473, 0.1976223, 0.2025083, 0.1971653, 0.2009866, 0.2022992, 
    0.2176784, 0.2228633, 0.2187544, 0.214001, 0.2185877, 0.2140497, 
    0.2061231, 0.2065106, 0.2014224, 0.2072845, 0.206794, 0.2046946, 
    0.2145764, 0.2025695, 0.1916149, 0.2092959, 0.1983277, 0.1910123, 
    0.1984383, 0.1941958, 0.193971, 0.2023256, 0.2020953, 0.1957219, 
    0.1837536, 0.1737093, 0.1683474, 0.1846378, 0.1777872, 0.1723011, 
    0.1912805, 0.1863299, 0.1861476, 0.1910618, 0.189579, 0.1911637, 
    0.1660194, 0.1663002, 0.1632531, 0.1726962, 0.1692982, 0.1692332, 
    0.1866185, 0.185738, 0.183803, 0.1944554, 0.1878936, 0.1843572, 
    0.1645128, 0.1611739, 0.1654865, 0.1674676, 0.1732864, 0.1793182, 
    0.1782852, 0.1799644, 0.1806711, 0.1824575, 0.1812101, 0.1796821, 
    0.1727975, 0.1810001, 0.1790856, 0.1820909, 0.1839266, 0.1824702, 
    0.1802306, 0.1785491, 0.1783706, 0.1801679, 0.1798219, 0.1800515, 
    0.1782534, 0.1707326, 0.165179, 0.1780285, 0.1716749,
  0.2328141, 0.2253507, 0.2235527, 0.2561473, 0.2486514, 0.2459111, 0.280061, 
    0.2749005, 0.2761213, 0.3008731, 0.2998164, 0.2962229, 0.2184264, 
    0.2138063, 0.209667, 0.2384951, 0.2267841, 0.2254802, 0.2729947, 
    0.2731359, 0.2619722, 0.2914295, 0.2903389, 0.2793564, 0.206498, 
    0.2038189, 0.2029108, 0.2194337, 0.2103137, 0.2083619, 0.2561122, 
    0.2471438, 0.2428971, 0.2763221, 0.2657825, 0.2653511, 0.1990098, 
    0.1978013, 0.1951801, 0.2082962, 0.1985353, 0.1937048, 0.2407465, 
    0.2322109, 0.2296394, 0.2653607, 0.2673402, 0.2678256, 0.1939786, 
    0.187762, 0.1823819, 0.1911756, 0.1887725, 0.1853522, 0.2262627, 
    0.225146, 0.2273801, 0.2677045, 0.2643768, 0.2698668, 0.1837924, 
    0.1829629, 0.1794883, 0.1842971, 0.182448, 0.1830351, 0.2240176, 
    0.225499, 0.2245524, 0.2692265, 0.2637211, 0.2574579, 0.1825373, 
    0.1837556, 0.1818831, 0.1876919, 0.1920198, 0.1933108, 0.2221532, 
    0.2253574, 0.2200859, 0.2534838, 0.248567, 0.2446133, 0.1823702, 
    0.1832367, 0.1770775, 0.197365, 0.1954164, 0.1967893, 0.2205968, 
    0.2237628, 0.2201617, 0.24115, 0.2416659, 0.2385316, 0.1788117, 
    0.1795344, 0.175938, 0.1973906, 0.1963828,
  0.204444, 0.2072698, 0.2067574, 0.2176633, 0.2135747, 0.2178392, 0.2335735, 
    0.2299278, 0.2262418, 0.2236743, 0.2212161, 0.2159656, 0.2084925, 
    0.2021631, 0.2008516, 0.2226151, 0.2189734, 0.2158672, 0.2217481, 
    0.2190054, 0.2204123, 0.2130173, 0.2136159, 0.2142838, 0.2027153, 
    0.206304, 0.2081103, 0.2174216, 0.2124261, 0.2099107, 0.2184698, 
    0.2157317, 0.2140991, 0.219043, 0.2140676, 0.2128523, 0.2107146, 
    0.2122156, 0.2090498, 0.2133374, 0.2115416, 0.2058555, 0.2109797, 
    0.2048368, 0.2043152, 0.2105579, 0.2080344, 0.2062403, 0.2067657, 
    0.2013219, 0.200346, 0.2065167, 0.2008361, 0.1984873, 0.2001425, 
    0.2000109, 0.1979567, 0.2059634, 0.2031755, 0.2030543, 0.1996704, 
    0.1920203, 0.1821725, 0.1973005, 0.1906978, 0.1843055, 0.197426, 
    0.1928427, 0.1902122, 0.2033072, 0.2016314, 0.1979146, 0.1774764, 
    0.1716716, 0.1653709, 0.1831256, 0.1775313, 0.1754184, 0.1897976, 
    0.186005, 0.1863624, 0.1977658, 0.1952214, 0.1950417, 0.1671808, 
    0.1680032, 0.1682307, 0.1742246, 0.1789841, 0.1745003, 0.1895942, 
    0.18645, 0.1821378, 0.1953169, 0.1920279, 0.1882636, 0.1707138, 
    0.1733059, 0.1777821, 0.1737445, 0.1800582,
  0.1874763, 0.1854456, 0.1814247, 0.1976035, 0.1998249, 0.1943721, 0.181789, 
    0.1794651, 0.1787239, 0.1732308, 0.1759064, 0.1783534, 0.1802338, 
    0.1753629, 0.1733582, 0.1895151, 0.1836687, 0.1836294, 0.1798311, 
    0.1776651, 0.1788806, 0.1808146, 0.1874484, 0.1917937, 0.1724441, 
    0.175578, 0.1767362, 0.1828668, 0.1839954, 0.1871086, 0.1845045, 
    0.1909551, 0.1983147, 0.195524, 0.2031294, 0.2073578, 0.1791757, 
    0.1824039, 0.1865295, 0.1908334, 0.1931793, 0.1944435, 0.2044816, 
    0.2137128, 0.2177168, 0.2139698, 0.2200673, 0.2263955, 0.1917258, 
    0.1921584, 0.1917933, 0.2003127, 0.2016572, 0.2016441, 0.2196665, 
    0.2220605, 0.2207931, 0.2291016, 0.2282213, 0.2269297, 0.1951355, 
    0.1926471, 0.1904399, 0.2039793, 0.2054035, 0.2021953, 0.226084, 
    0.2211898, 0.2169362, 0.2291686, 0.2223285, 0.2205108, 0.192067, 
    0.1860932, 0.1825772, 0.1986128, 0.19397, 0.1925947, 0.2149823, 
    0.2083118, 0.2072918, 0.2146216, 0.2106358, 0.2068996, 0.1826895, 
    0.1812841, 0.1783689, 0.1925931, 0.1915429, 0.1877338, 0.2053726, 
    0.2062912, 0.2117327, 0.2081459, 0.2069673, 0.2057144, 0.1760216, 
    0.1741731, 0.1701998, 0.1882237, 0.187264,
  0.1639496, 0.1595451, 0.156531, 0.1652171, 0.1610244, 0.1591977, 0.1557436, 
    0.1509242, 0.147754, 0.145687, 0.1427514, 0.1401382, 0.155261, 0.1537484, 
    0.1506867, 0.1573244, 0.1542185, 0.1504657, 0.1449548, 0.139431, 
    0.1368212, 0.1376683, 0.1318312, 0.1290433, 0.1428579, 0.1331931, 
    0.1306754, 0.1459978, 0.1365148, 0.1328484, 0.1346847, 0.129936, 
    0.1305152, 0.1280837, 0.1281873, 0.1286501, 0.1295359, 0.1266263, 
    0.12501, 0.1320954, 0.1341981, 0.1366763, 0.1332892, 0.141581, 0.1454187, 
    0.1322034, 0.1391025, 0.1443336, 0.1230571, 0.1240539, 0.1252189, 
    0.1361701, 0.1384341, 0.1381979, 0.1478914, 0.1534673, 0.1557051, 
    0.1472054, 0.1534983, 0.1586755, 0.1258428, 0.131171, 0.1332238, 
    0.1397339, 0.1444615, 0.1440398, 0.1596013, 0.1657794, 0.167528, 0.16337, 
    0.1698887, 0.1687638, 0.1377382, 0.146675, 0.1497508, 0.1477413, 
    0.155737, 0.1595023, 0.1687649, 0.1701479, 0.1669537, 0.1701636, 
    0.1695872, 0.1655654, 0.1530678, 0.1561455, 0.1565032, 0.1594906, 
    0.1585625, 0.1550934, 0.1625452, 0.1582287, 0.1546297, 0.1649762, 
    0.1584144, 0.1544651, 0.1558895, 0.1566933, 0.156946, 0.1553478, 0.1537159,
  0.1353782, 0.1312087, 0.1292458, 0.1426762, 0.1361229, 0.1328902, 
    0.1535928, 0.1433089, 0.1388196, 0.1573098, 0.146523, 0.1389918, 
    0.1245651, 0.1150763, 0.109313, 0.1279398, 0.1192965, 0.1135766, 
    0.1309429, 0.1231705, 0.1198923, 0.1323208, 0.1258093, 0.1217002, 
    0.1040016, 0.1016777, 0.09872911, 0.1067144, 0.1047865, 0.1015466, 
    0.1154291, 0.1124931, 0.1088241, 0.1172297, 0.1116155, 0.1078881, 
    0.09788425, 0.09889922, 0.0999926, 0.09980367, 0.1035499, 0.1045499, 
    0.1056143, 0.1055134, 0.1063924, 0.1026411, 0.1048483, 0.107031, 
    0.1008385, 0.09706043, 0.09352417, 0.1052834, 0.09941827, 0.09489581, 
    0.1068266, 0.1028343, 0.09999228, 0.1077049, 0.1068426, 0.1064215, 
    0.08877205, 0.08181074, 0.08057696, 0.09097475, 0.08514158, 0.08170754, 
    0.09858683, 0.09541271, 0.09283178, 0.1056114, 0.09951932, 0.09540126, 
    0.07911389, 0.07714377, 0.07695907, 0.08063359, 0.07975329, 0.08066572, 
    0.09082519, 0.08779536, 0.08894471, 0.09267303, 0.09253707, 0.09651057, 
    0.07706194, 0.0776449, 0.07805382, 0.08135448, 0.08540493, 0.08491925, 
    0.09154148, 0.09411108, 0.09483948, 0.09866248, 0.1024592, 0.1038351, 
    0.07768513, 0.07748754, 0.07787821, 0.08415257, 0.08371783,
  0.1382949, 0.1450226, 0.148034, 0.1351843, 0.1423517, 0.1455969, 0.1269834, 
    0.1332947, 0.1362588, 0.1188061, 0.1254395, 0.128265, 0.1504975, 
    0.1513442, 0.1490947, 0.148807, 0.149872, 0.1480099, 0.1397791, 
    0.1434865, 0.1443396, 0.1318148, 0.1365135, 0.1382835, 0.1487013, 
    0.1486881, 0.1485823, 0.146389, 0.1456712, 0.1477453, 0.1452807, 
    0.1472689, 0.1519227, 0.1412855, 0.1469412, 0.151781, 0.1509573, 
    0.1542943, 0.1552909, 0.1527777, 0.1558307, 0.1582843, 0.154592, 
    0.1606407, 0.1639641, 0.1554668, 0.1610759, 0.1626997, 0.1541734, 
    0.1541477, 0.1518399, 0.1604304, 0.1583867, 0.1580848, 0.1672571, 
    0.1651968, 0.1613963, 0.1653595, 0.1633147, 0.1615627, 0.1508166, 
    0.1512521, 0.1531667, 0.1548624, 0.1537739, 0.1559115, 0.1594255, 
    0.1581944, 0.1571706, 0.1596704, 0.1558136, 0.156253, 0.1532934, 
    0.1551352, 0.156336, 0.1558671, 0.1586895, 0.160724, 0.158261, 0.158468, 
    0.1603837, 0.1562793, 0.1582433, 0.1591779, 0.1579367, 0.1617875, 
    0.1627547, 0.1620818, 0.1650384, 0.1638088, 0.1614345, 0.1611486, 
    0.1601361, 0.1606927, 0.1607834, 0.1580767, 0.1616362, 0.1614227, 
    0.1611511, 0.1609218, 0.158991,
  0.1428538, 0.1445044, 0.1425923, 0.1426579, 0.1413944, 0.1407125, 
    0.1364104, 0.1366594, 0.1363738, 0.132962, 0.1319296, 0.1338147, 
    0.1429807, 0.1430847, 0.1434638, 0.1399993, 0.1414684, 0.1439629, 
    0.1383283, 0.1417851, 0.1464691, 0.1367006, 0.1418087, 0.1424577, 
    0.1437016, 0.145293, 0.1442515, 0.1449031, 0.1476569, 0.1505536, 
    0.1447543, 0.1483661, 0.1524974, 0.1446298, 0.1466715, 0.147372, 
    0.1469412, 0.1494225, 0.1517926, 0.1527238, 0.156586, 0.158306, 
    0.1534151, 0.1582753, 0.1619965, 0.1515539, 0.1578692, 0.1613436, 
    0.1536035, 0.1559664, 0.1576068, 0.1609645, 0.1624408, 0.166122, 
    0.1647256, 0.1710236, 0.174675, 0.1640714, 0.1686623, 0.1714816, 
    0.158515, 0.162247, 0.1654732, 0.1683774, 0.1704258, 0.1733287, 
    0.1775742, 0.1817226, 0.1841532, 0.1710595, 0.1750595, 0.1757429, 
    0.1682188, 0.173983, 0.1759125, 0.1771324, 0.1809456, 0.1844898, 0.18458, 
    0.1847741, 0.1817765, 0.1773918, 0.1762646, 0.1798744, 0.1793412, 
    0.1851471, 0.1884616, 0.1861663, 0.1875532, 0.1855837, 0.1784803, 
    0.1789475, 0.1800691, 0.1757767, 0.1791561, 0.1790625, 0.1870868, 
    0.1856772, 0.1812662, 0.1849439, 0.1827552,
  0.1114668, 0.1117572, 0.1137109, 0.1123473, 0.1090506, 0.1091674, 
    0.1066714, 0.1048104, 0.1053871, 0.1061258, 0.1047961, 0.1042288, 
    0.1143955, 0.1188063, 0.1245094, 0.1099888, 0.116806, 0.1214506, 
    0.1079257, 0.1128635, 0.1143611, 0.1051767, 0.1077919, 0.110173, 
    0.1251327, 0.1245165, 0.1238515, 0.1247278, 0.1264436, 0.1277844, 
    0.1194365, 0.1244638, 0.1256402, 0.1139666, 0.1197496, 0.119506, 
    0.1252479, 0.1245234, 0.1231315, 0.1282175, 0.1265963, 0.1276615, 
    0.1240689, 0.1243562, 0.1256312, 0.1186379, 0.1200207, 0.1232827, 
    0.1222743, 0.1204777, 0.119525, 0.1248277, 0.1259445, 0.1263142, 
    0.1279189, 0.1308628, 0.1350332, 0.1256219, 0.1326889, 0.1359928, 
    0.1201318, 0.1232656, 0.1298773, 0.1284368, 0.132803, 0.1360237, 
    0.1384837, 0.1423043, 0.1415664, 0.1382871, 0.1405343, 0.1397824, 
    0.131799, 0.1329814, 0.1332365, 0.1354107, 0.1343369, 0.1333424, 
    0.1415186, 0.1380852, 0.1352166, 0.1379745, 0.1361696, 0.1341835, 
    0.1328081, 0.1331753, 0.1347166, 0.1341383, 0.1334959, 0.1333819, 
    0.1316389, 0.1315629, 0.1319548, 0.1327208, 0.1304544, 0.1307182, 
    0.1372361, 0.1406366, 0.1418632, 0.1364852, 0.1397609,
  0.1602387, 0.1568671, 0.1544906, 0.1440604, 0.1443709, 0.1444191, 
    0.1284406, 0.1277434, 0.1277922, 0.128046, 0.1280519, 0.1289813, 
    0.1534733, 0.150717, 0.1503597, 0.1430183, 0.140761, 0.1419737, 
    0.1285734, 0.1308771, 0.1329144, 0.1288784, 0.1297022, 0.130541, 
    0.1495953, 0.1486224, 0.1488258, 0.1436143, 0.1437625, 0.1431728, 
    0.1346518, 0.1323624, 0.1311874, 0.1310046, 0.1309152, 0.1293972, 
    0.1491942, 0.1499555, 0.1462928, 0.1411681, 0.1367763, 0.1327885, 
    0.1286456, 0.1237259, 0.1212917, 0.1249014, 0.1192282, 0.1162069, 
    0.1431972, 0.1392267, 0.1355784, 0.1299733, 0.1258703, 0.1229684, 
    0.1187575, 0.1165072, 0.1165477, 0.1147363, 0.1145243, 0.1140298, 
    0.1292798, 0.1212466, 0.1181903, 0.1211085, 0.1172793, 0.1165111, 
    0.1171926, 0.12089, 0.1232592, 0.1144994, 0.1198958, 0.1221344, 
    0.1154956, 0.1157786, 0.1169998, 0.1167669, 0.1212647, 0.1224213, 
    0.1242012, 0.1284865, 0.1284122, 0.121344, 0.1229231, 0.1232181, 
    0.1210874, 0.1234303, 0.1256993, 0.125475, 0.1273831, 0.1284126, 
    0.1291642, 0.1268377, 0.1245345, 0.1226114, 0.1213361, 0.119859, 
    0.1271431, 0.1290349, 0.1276836, 0.1264341, 0.1261583,
  0.1050755, 0.1062234, 0.1061448, 0.1020185, 0.1024253, 0.1032896, 
    0.1002943, 0.1006925, 0.09957704, 0.1066907, 0.1065698, 0.1051571, 
    0.1051281, 0.102196, 0.1024118, 0.1017433, 0.0991314, 0.09848049, 
    0.09843103, 0.09766504, 0.097927, 0.1028765, 0.1005712, 0.09923952, 
    0.1022633, 0.1039979, 0.1044579, 0.09935891, 0.1015145, 0.1021418, 
    0.0987502, 0.1016327, 0.1025257, 0.09918553, 0.1010293, 0.1031687, 
    0.1070372, 0.1116234, 0.1150643, 0.1051012, 0.1092137, 0.1112501, 
    0.1051245, 0.1050213, 0.1061022, 0.1046324, 0.1060196, 0.1071381, 
    0.120111, 0.1264709, 0.1298779, 0.1138941, 0.1209193, 0.1252851, 
    0.107301, 0.1093941, 0.11171, 0.1071246, 0.1096588, 0.1118321, 0.1347528, 
    0.1393142, 0.1410836, 0.127227, 0.1311932, 0.1327865, 0.114323, 
    0.1208021, 0.1235724, 0.1144281, 0.1190242, 0.1206391, 0.1444131, 
    0.145172, 0.1450475, 0.1341155, 0.1370124, 0.1383893, 0.1265653, 
    0.1283886, 0.1298017, 0.1235624, 0.1282434, 0.1312317, 0.1427317, 
    0.1436867, 0.1469251, 0.1394262, 0.1414875, 0.1459295, 0.1314368, 
    0.1366657, 0.1385289, 0.1311646, 0.1338378, 0.1359334, 0.1485552, 
    0.1532829, 0.1562486, 0.1476973, 0.1523531,
  0.1915207, 0.1905512, 0.1891114, 0.1900187, 0.1928829, 0.1920616, 
    0.1788477, 0.1781291, 0.1769752, 0.1696773, 0.169655, 0.1701644, 
    0.187976, 0.1816119, 0.1834482, 0.192444, 0.1906275, 0.1885915, 
    0.1794916, 0.1827076, 0.1870105, 0.1739968, 0.1799391, 0.1853353, 
    0.1876314, 0.1864454, 0.1837543, 0.1892748, 0.1923203, 0.1959099, 
    0.1907911, 0.1988162, 0.2028057, 0.191971, 0.199615, 0.2028668, 0.184936, 
    0.1882321, 0.1896854, 0.1986764, 0.2011138, 0.2025274, 0.2051796, 
    0.203412, 0.2006076, 0.1991198, 0.2001319, 0.1999938, 0.1910143, 
    0.192018, 0.1954547, 0.2032, 0.2045579, 0.2040587, 0.2031571, 0.2026904, 
    0.2030691, 0.198571, 0.2013117, 0.2038108, 0.1976015, 0.2067915, 
    0.2086159, 0.2026002, 0.2071473, 0.2082788, 0.2025556, 0.2026761, 
    0.1998926, 0.2030682, 0.2004396, 0.1965656, 0.2099271, 0.2168364, 
    0.2195687, 0.2093928, 0.2117628, 0.2133301, 0.1996985, 0.197555, 
    0.1922587, 0.1934512, 0.192504, 0.1924015, 0.2211165, 0.2104659, 
    0.2051557, 0.2137458, 0.205901, 0.2018786, 0.1900305, 0.1892061, 
    0.1922204, 0.1943211, 0.2013324, 0.2001679, 0.2019928, 0.1955626, 
    0.1910436, 0.1977003, 0.1956208,
  0.1786886, 0.1833761, 0.182936, 0.167746, 0.1711043, 0.1717877, 0.1562743, 
    0.1560527, 0.1590466, 0.1480945, 0.1545533, 0.1568717, 0.1813385, 
    0.1727088, 0.1717167, 0.1711712, 0.1689125, 0.165551, 0.1609344, 
    0.1642672, 0.1635927, 0.1605262, 0.1660524, 0.1657453, 0.1678452, 
    0.1642451, 0.1616925, 0.1640777, 0.1643642, 0.1623019, 0.163319, 
    0.1677254, 0.1734749, 0.1641901, 0.1677097, 0.1693747, 0.1598094, 
    0.1555314, 0.1559358, 0.1617846, 0.1613723, 0.1613546, 0.1744929, 
    0.1762118, 0.1798715, 0.1715388, 0.1774809, 0.1809742, 0.1538051, 
    0.1546992, 0.1531337, 0.1675038, 0.1709409, 0.170484, 0.1796484, 
    0.1820846, 0.1844894, 0.1858571, 0.1907896, 0.1913448, 0.1550318, 
    0.1598441, 0.156537, 0.1721136, 0.1702973, 0.1705465, 0.1889088, 
    0.181659, 0.1813747, 0.1922163, 0.1849335, 0.1813839, 0.1604174, 
    0.1618205, 0.162083, 0.1688964, 0.1680832, 0.1637787, 0.1786449, 
    0.1716461, 0.16596, 0.1759826, 0.1694941, 0.1653446, 0.1609978, 
    0.1657248, 0.1669308, 0.1632226, 0.1610157, 0.1619247, 0.1615189, 
    0.1582473, 0.1569887, 0.1638287, 0.1625439, 0.1635265, 0.1712507, 
    0.179959, 0.1799442, 0.1672631, 0.1770737,
  0.2190626, 0.2161675, 0.2124575, 0.2151826, 0.2086686, 0.2061593, 
    0.2064152, 0.2034399, 0.1979037, 0.2011914, 0.192725, 0.1907427, 
    0.206601, 0.2032417, 0.2026785, 0.2008825, 0.1951693, 0.1938006, 
    0.1935272, 0.1936183, 0.1935009, 0.1886067, 0.190855, 0.1953703, 
    0.2006611, 0.1967442, 0.1991313, 0.1929758, 0.1959505, 0.1954374, 
    0.1948512, 0.203792, 0.2057316, 0.1947606, 0.2063612, 0.2107576, 
    0.2026935, 0.2014569, 0.2010473, 0.1977097, 0.1999278, 0.1992519, 
    0.2057605, 0.2057374, 0.2046032, 0.2137366, 0.2117251, 0.2107314, 
    0.1978284, 0.1996669, 0.2012285, 0.202851, 0.2026321, 0.2026318, 
    0.2057471, 0.2081716, 0.2079574, 0.2091661, 0.2094062, 0.2091158, 
    0.1973222, 0.1981285, 0.1977272, 0.2027561, 0.2015419, 0.1968763, 
    0.2093275, 0.2066158, 0.2043409, 0.2050741, 0.2039009, 0.2029746, 
    0.1941545, 0.190312, 0.1831876, 0.1987242, 0.1962608, 0.1952614, 
    0.2027334, 0.1972917, 0.2024268, 0.2021926, 0.1986063, 0.2034607, 
    0.181661, 0.1801108, 0.1811988, 0.1904286, 0.1912836, 0.1912515, 
    0.2080938, 0.2137125, 0.224667, 0.2090217, 0.2226768, 0.2244089, 
    0.1799948, 0.1855928, 0.1905904, 0.1959832, 0.2028412,
  0.2363871, 0.2310137, 0.2275852, 0.2397519, 0.2378715, 0.2391831, 0.270887, 
    0.2670993, 0.2654123, 0.2675422, 0.2742962, 0.2755051, 0.2293099, 
    0.233057, 0.2325758, 0.2442331, 0.247789, 0.2447284, 0.2689262, 
    0.2779264, 0.2778774, 0.2780661, 0.2794837, 0.2799218, 0.2292865, 
    0.223557, 0.2233916, 0.2446221, 0.2425748, 0.2424671, 0.2795719, 
    0.2866049, 0.2844692, 0.2829563, 0.2805229, 0.2772895, 0.228307, 
    0.2256315, 0.2290545, 0.2481035, 0.2468491, 0.2458177, 0.2804992, 
    0.2848791, 0.2817129, 0.2751534, 0.2799759, 0.2863012, 0.2313857, 
    0.2375565, 0.2440142, 0.2485435, 0.2558631, 0.2578455, 0.2849799, 
    0.2769746, 0.273105, 0.2868959, 0.2846403, 0.2828279, 0.2495223, 
    0.255291, 0.2502186, 0.2611667, 0.2678204, 0.2652672, 0.2677513, 
    0.2659397, 0.2641079, 0.2783761, 0.2705274, 0.2651047, 0.2500214, 
    0.2407222, 0.2320614, 0.2642207, 0.2563878, 0.2503784, 0.2596502, 
    0.2562346, 0.2570219, 0.2645656, 0.2599223, 0.255474, 0.2288296, 
    0.2171425, 0.2138653, 0.2479661, 0.2364154, 0.2348483, 0.2546183, 
    0.2554798, 0.2620098, 0.2596889, 0.2651418, 0.2680561, 0.2138027, 
    0.2154066, 0.2126942, 0.2365976, 0.2433262,
  0.2273601, 0.2264391, 0.2249806, 0.2255498, 0.2239716, 0.225776, 0.2341366, 
    0.2271899, 0.2237888, 0.2365928, 0.2294157, 0.2291263, 0.2244227, 
    0.2252293, 0.2251894, 0.2243496, 0.2264393, 0.2273743, 0.2253674, 
    0.224435, 0.226916, 0.2306219, 0.2329614, 0.2306426, 0.2281481, 
    0.2254229, 0.2233813, 0.2320441, 0.2302232, 0.2302986, 0.2316897, 
    0.2338728, 0.237324, 0.2318275, 0.2308813, 0.2316375, 0.2269405, 
    0.2279114, 0.2335363, 0.2294652, 0.2329853, 0.2355096, 0.237585, 
    0.2372299, 0.2394412, 0.2318557, 0.2359824, 0.2397066, 0.2362248, 
    0.2384186, 0.2411703, 0.2406262, 0.2446066, 0.2434119, 0.2428299, 
    0.2489082, 0.2499716, 0.2461069, 0.2535728, 0.2554342, 0.2422964, 
    0.2410934, 0.2357847, 0.2438002, 0.246578, 0.2471658, 0.2526763, 
    0.2536096, 0.2476416, 0.2481783, 0.2420948, 0.2422484, 0.2351049, 
    0.2339057, 0.2263373, 0.2454067, 0.2410341, 0.2382855, 0.2404874, 
    0.2374443, 0.2392842, 0.239357, 0.2421721, 0.2457046, 0.2251948, 
    0.2222316, 0.2207261, 0.2368596, 0.2343885, 0.2265344, 0.2401103, 
    0.2402156, 0.2356424, 0.2496521, 0.2496633, 0.2449977, 0.2161435, 
    0.211295, 0.2062158, 0.2196096, 0.217275,
  0.1833392, 0.1814924, 0.1803719, 0.1779939, 0.1768701, 0.176074, 0.1634538, 
    0.1678145, 0.1710857, 0.1644397, 0.1675935, 0.1695061, 0.1830664, 
    0.1833141, 0.1823932, 0.1813454, 0.1878084, 0.1877795, 0.1772014, 
    0.1823444, 0.1833619, 0.1713593, 0.1746094, 0.1751955, 0.1816076, 
    0.1776618, 0.1789077, 0.1878611, 0.1857078, 0.1825854, 0.1847088, 
    0.1824234, 0.1797517, 0.1735295, 0.1732109, 0.1722764, 0.1811599, 
    0.180442, 0.178427, 0.1818759, 0.1808412, 0.1791587, 0.178409, 0.1767042, 
    0.1759668, 0.1732458, 0.1743387, 0.1759574, 0.1789876, 0.1809032, 
    0.1813175, 0.179189, 0.1849938, 0.1870098, 0.1775593, 0.183135, 
    0.1853722, 0.1773289, 0.1833863, 0.1853209, 0.184155, 0.18352, 0.1796999, 
    0.1892099, 0.1900401, 0.1876739, 0.1882673, 0.1859271, 0.1835845, 
    0.1846513, 0.1807886, 0.1759426, 0.1806132, 0.1761451, 0.1756252, 
    0.1861437, 0.1846994, 0.1806708, 0.1805478, 0.1782488, 0.1746423, 
    0.1748901, 0.1683411, 0.162845, 0.1711306, 0.1672867, 0.1652438, 
    0.1796088, 0.1778824, 0.1749175, 0.1725637, 0.1698459, 0.1680615, 
    0.1605286, 0.1572239, 0.1567249, 0.163386, 0.1595778, 0.1579816, 
    0.1756621, 0.1677156,
  0.1768353, 0.1704365, 0.1662122, 0.170723, 0.1668689, 0.1620558, 0.1627614, 
    0.1571805, 0.1536792, 0.1574781, 0.1557824, 0.151551, 0.1634641, 
    0.158519, 0.1565732, 0.1578867, 0.1537219, 0.1524752, 0.1521743, 
    0.1523545, 0.1517183, 0.1499506, 0.1510862, 0.1499685, 0.1531481, 
    0.1518757, 0.149415, 0.1521942, 0.1532604, 0.1532426, 0.1546461, 
    0.1554156, 0.1561447, 0.1512384, 0.1552559, 0.156931, 0.1491171, 
    0.1478736, 0.1456751, 0.1537527, 0.1523206, 0.1502036, 0.1552065, 
    0.1527256, 0.1532962, 0.1574454, 0.160001, 0.1599603, 0.1456407, 
    0.1426908, 0.139314, 0.1497785, 0.1473956, 0.1457293, 0.1549507, 
    0.1572608, 0.1574807, 0.1613142, 0.1583218, 0.1542286, 0.139235, 
    0.1382236, 0.1372044, 0.1475934, 0.1460287, 0.1456109, 0.1560339, 
    0.1503131, 0.1460616, 0.1498879, 0.1413872, 0.1363711, 0.1380679, 
    0.1366222, 0.1371197, 0.1445503, 0.1424511, 0.1413202, 0.1424686, 
    0.1437623, 0.1440656, 0.1349784, 0.1398705, 0.1434058, 0.138155, 
    0.1375185, 0.1402052, 0.1415428, 0.1436862, 0.1436375, 0.144942, 
    0.1449981, 0.1463917, 0.1430753, 0.1459787, 0.150064, 0.1418546, 
    0.1447684, 0.1497619, 0.1454354, 0.149112,
  0.1233806, 0.1299262, 0.1329367, 0.1281853, 0.1356412, 0.1379512, 
    0.1329578, 0.1425893, 0.1468584, 0.1334201, 0.1453158, 0.1492854, 
    0.1328756, 0.1306882, 0.1301605, 0.1370767, 0.1355338, 0.1321272, 
    0.1446117, 0.1415721, 0.1392124, 0.1503075, 0.1456869, 0.143813, 
    0.1303605, 0.1271376, 0.1209919, 0.1317295, 0.1305591, 0.1253362, 
    0.1381487, 0.1354873, 0.1300382, 0.1400403, 0.1343057, 0.1309104, 
    0.1169696, 0.1072834, 0.1040777, 0.1214785, 0.1125156, 0.1067991, 
    0.1209835, 0.1080683, 0.1026791, 0.1213782, 0.1082171, 0.1063813, 
    0.1044694, 0.09722704, 0.0961274, 0.1016289, 0.09655076, 0.09794204, 
    0.1007176, 0.1026715, 0.1038659, 0.1067826, 0.1079552, 0.1073005, 
    0.09593774, 0.09795097, 0.09939069, 0.1004332, 0.1028993, 0.1029212, 
    0.1028891, 0.1009039, 0.09836306, 0.1023176, 0.09687418, 0.09234102, 
    0.09733045, 0.09784158, 0.09686849, 0.1021902, 0.1000225, 0.09701466, 
    0.09519687, 0.08951161, 0.08669902, 0.088146, 0.08186313, 0.07960083, 
    0.09664916, 0.09513067, 0.09237097, 0.0942224, 0.0887329, 0.0881855, 
    0.08329523, 0.08116913, 0.08005256, 0.07773824, 0.07640599, 0.07517501, 
    0.0910221, 0.08911258, 0.08775266, 0.08715925, 0.08547039,
  0.1688406, 0.1710348, 0.171356, 0.1672868, 0.1718615, 0.1727286, 0.1633426, 
    0.1644738, 0.1644144, 0.1661194, 0.1670091, 0.1660045, 0.1718054, 
    0.1682719, 0.1654034, 0.1748282, 0.1699753, 0.1676045, 0.1658645, 
    0.1670622, 0.1647154, 0.1662265, 0.1661081, 0.165916, 0.1615234, 
    0.1551331, 0.1514707, 0.1645463, 0.1607642, 0.1564291, 0.1634826, 
    0.1587933, 0.1555076, 0.1627442, 0.158357, 0.155075, 0.1489802, 
    0.1424965, 0.1399803, 0.1511063, 0.1454895, 0.1420271, 0.1513158, 
    0.1447111, 0.1437266, 0.1521958, 0.1472662, 0.1482003, 0.1372176, 
    0.1331309, 0.1292118, 0.1412891, 0.1362127, 0.1305578, 0.1437601, 
    0.1430719, 0.1433737, 0.150409, 0.1526376, 0.1560405, 0.1252463, 
    0.1210408, 0.1199998, 0.1261948, 0.123648, 0.1241905, 0.1430184, 
    0.1435985, 0.1426001, 0.1581886, 0.1569205, 0.15503, 0.1197255, 
    0.1180008, 0.1192861, 0.126414, 0.1271208, 0.1281044, 0.1430035, 
    0.1451576, 0.1436733, 0.1498344, 0.1410937, 0.1336634, 0.1188039, 
    0.1202592, 0.1214578, 0.1255444, 0.1264641, 0.1251924, 0.1382788, 
    0.125625, 0.1243998, 0.1295239, 0.126437, 0.1259565, 0.1198862, 
    0.1209796, 0.1250039, 0.1273838, 0.1288886 ;

 area = 0.000138535035537854, 0.000138063242676441, 5.51133351740581e-05, 
    0.000350351563033784, 0.000349283468177034, 0.000139459179024405, 
    0.000356644999159883, 0.000355762606968429, 0.000142093741826655, 
    0.000144164429551706, 0.000143858593374666, 5.74698205985682e-05, 
    0.000137512973925224, 0.00013709691415187, 5.47414700454348e-05, 
    0.000348032852535342, 0.000347084025582322, 0.000138611239906833, 
    0.000354720920990366, 0.000353924965687112, 0.000141382596205829, 
    0.000143495040191689, 0.000143215599555958, 5.72202057728467e-05, 
    0.000136621526727059, 0.000136270294293906, 5.44275208617861e-05, 
    0.000345996716970601, 0.000345191311810852, 0.000137891406276323, 
    0.000353007300225509, 0.000352323972686935, 0.0001407720046366, 
    0.000142891821216884, 0.000142649689936032, 5.70038865267309e-05, 
    0.000135879563900365, 0.000135599984935344, 5.41776043392406e-05, 
    0.000344293376801085, 0.000343649664097871, 0.000137316047087783, 
    0.000351558750150899, 0.000351008077914795, 0.000140279905662028, 
    0.000142377566253734, 0.000142181139436531, 5.68283813074782e-05, 
    0.000135301131646374, 0.000135098141809231, 5.39961435185002e-05, 
    0.000342960495355738, 0.000342491775166504, 0.000136897078836035, 
    0.000350416658918027, 0.00035001335752274, 0.00013991948065301, 
    0.000141969647815823, 0.000141825125025086, 5.66992425861007e-05, 
    0.000134896237903517, 0.000134773166429464, 5.38861220302414e-05, 
    0.00034202508027183, 0.000341740372763005, 0.000136642583755051, 
    0.000349610968386061, 0.000349365092423242, 0.000139699736350274, 
    0.000141680693775172, 0.000141592327806752, 5.66202794187052e-05, 
    0.000134671432986883, 0.000134630200066165, 5.3849260799652e-05, 
    0.000341504897264425, 0.000341409424936482, 0.000136557241461346, 
    0.000349161509538827, 0.000349078910701538, 0.00013962591475864, 
    0.000141519098339092, 0.000141489371108393, 5.65937148161597e-05, 
    0.000134630200066165, 0.000134671432986883, 5.38861220302414e-05, 
    0.000341409424936482, 0.000341504897264425, 0.000136642583755051, 
    0.000349078910701538, 0.000349161509538827, 0.000139699736350274, 
    0.000141489371108393, 0.000141519098339092, 5.66202794187052e-05, 
    0.000134773166429464, 0.000134896237903517, 5.39961435185002e-05, 
    0.000341740372763005, 0.00034202508027183 ;

 lat = -43.1880092162786, -43.4251557914009, -43.5630005995731, 
    -42.3612436665401, -42.5978863344025, -42.7354642114613, 
    -41.0266990661296, -41.2621122848379, -41.399016975171, 
    -40.2038645450768, -40.4382645514851, -40.5746054270778, 
    -43.6942519279646, -43.8927912645738, -44.0070271956363, 
    -42.8664791346531, -43.0646938085549, -43.1787609186728, 
    -41.5294192763691, -41.7267599148945, -41.8403528927482, 
    -40.7044880945559, -40.9010746810136, -41.0142512786351, 
    -44.1148510165636, -44.2758447890606, -44.3670849826627, 
    -43.286437451671, -43.4472331078255, -43.5383726205395, 
    -41.9476012104333, -42.1077924196086, -42.1986079661906, 
    -41.1211183292902, -41.2807615219073, -41.3712778144978, 
    -44.4520614974551, -44.5763786122228, -44.6451168488014, 
    -43.6232629149409, -43.7474670128113, -43.8161494525006, 
    -42.2832086436371, -42.4070101005765, -42.4754806567305, 
    -41.4556071611961, -41.5790245116986, -41.6472892415569, 
    -44.7077067917174, -44.7960227295218, -44.842633221219, 
    -43.8786927360161, -43.9669495608533, -44.0135320282192, 
    -42.5378376701362, -42.625842470155, -42.6722970285562, 
    -41.7094629044609, -41.7972155906693, -41.8435402072463, 
    -44.8831777701286, -44.9359746369799, -44.960712147569, 
    -44.0540539833997, -44.1068239163782, -44.1315497755592, 
    -42.7127105890533, -42.765343372397, -42.7900065290456, 
    -41.8838424889767, -41.9363328110146, -41.9609301708143, 
    -44.9794330895693, -44.9969999412459, -45, -44.1502623106946, 
    -44.1678215955947, -44.1708203932499, -42.8086722728506, 
    -42.8261881688884, -42.8291796067501, -41.9795465246935, 
    -41.9970163922116, -42, -44.9969999412459, -44.9794330895693, 
    -44.960712147569, -44.1678215955947, -44.1502623106946, 
    -44.1315497755592, -42.8261881688884, -42.8086722728506, 
    -42.7900065290456, -41.9970163922116, -41.9795465246935, 
    -41.9609301708143, -44.9359746369799, -44.8831777701286, 
    -44.842633221219, -44.1068239163782, -44.0540539833997 ;

 lon = 339.82917960675, 341.17082039325, 342, 339.82917960675, 
    341.17082039325, 342, 339.82917960675, 341.17082039325, 342, 
    339.82917960675, 341.17082039325, 342, 342.82917960675, 344.17082039325, 
    345, 342.82917960675, 344.17082039325, 345, 342.82917960675, 
    344.17082039325, 345, 342.82917960675, 344.17082039325, 345, 
    345.82917960675, 347.17082039325, 348, 345.82917960675, 347.17082039325, 
    348, 345.82917960675, 347.17082039325, 348, 345.82917960675, 
    347.17082039325, 348, 348.82917960675, 350.17082039325, 351, 
    348.82917960675, 350.17082039325, 351, 348.82917960675, 350.17082039325, 
    351, 348.82917960675, 350.17082039325, 351, 351.82917960675, 
    353.17082039325, 354, 351.82917960675, 353.17082039325, 354, 
    351.82917960675, 353.17082039325, 354, 351.82917960675, 353.17082039325, 
    354, 354.82917960675, 356.17082039325, 357, 354.82917960675, 
    356.17082039325, 357, 354.82917960675, 356.17082039325, 357, 
    354.82917960675, 356.17082039325, 357, 357.82917960675, 359.17082039325, 
    360, 357.82917960675, 359.17082039325, 360, 357.82917960675, 
    359.17082039325, 360, 357.82917960675, 359.17082039325, 360, 
    0.829179606750063, 2.17082039324994, 3, 0.829179606750063, 
    2.17082039324994, 3, 0.829179606750063, 2.17082039324994, 3, 
    0.829179606750063, 2.17082039324994, 3, 3.82917960675006, 
    5.17082039324993, 6, 3.82917960675006, 5.17082039324993 ;

 time = 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 396, 424, 
    455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 820, 850, 
    881, 911, 942, 973, 1003, 1034, 1064, 1095 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365,
  365, 396,
  396, 424,
  424, 455,
  455, 485,
  485, 516,
  516, 546,
  546, 577,
  577, 608,
  608, 638,
  638, 669,
  669, 699,
  699, 730,
  730, 761,
  761, 789,
  789, 820,
  820, 850,
  850, 881,
  881, 911,
  911, 942,
  942, 973,
  973, 1003,
  1003, 1034,
  1034, 1064,
  1064, 1095 ;
}
