// Purpose: CDL file to generate netCDF test file for NCO

// Usage:
// netCDF4: ncgen arguments depend on version:
// "-k netCDF-4" for netCDF >= 3.6.3, "-k hdf5" for netCDF < 3.6.3
// "-k netCDF-4 classic model" for netCDF >= 3.6.3, "-k hdf5-nc3" for netCDF < 3.6.3
// /usr/local/bin/ncgen -k netCDF-4 -b -o in_4.nc in.cdl
// /usr/local/bin/ncgen -k netCDF-4 -b -o ${HOME}/nco/data/in_4.nc ${HOME}/nco/data/in.cdl

// URL: 
// http://dust.ess.uci.edu/nco/in.nc
// http://dust.ess.uci.edu/nco/in_4.nc

// netCDF3:
// ncgen -b -o in.nc in.cdl
// ncgen -b -o ${HOME}/nco/data/in.nc ${HOME}/nco/data/in.cdl
// scp ~/nco/data/in.cdl esmf.ess.uci.edu:nco/data
// scp ~/nco/data/in.nc dust.ess.uci.edu:/var/www/html/nco
// scp ~/nco/data/in.nc dust.ess.uci.edu:/data/home/www/html/dodsdata
// mswrite -t 365 ~/nco/data/in.nc /ZENDER/tmp/in.nc
// mswrite -t 365 ~/nco/data/in.nc /ZENDER/tmp/h0001.nc
// mswrite -t 365 ~/nco/data/in.nc /ZENDER/tmp/h0002.nc
// mswrite -t 365 ~/nco/data/in.nc /ZENDER/tmp/h0003.nc
// mswrite -t 365 ~/nco/data/in.nc /ZENDER/tmp/h0004.nc
// msrcp -period 365 ~/nco/data/in.nc mss:/ZENDER/tmp/in.nc
// msrcp -period 365 ~/nco/data/in.nc mss:/ZENDER/tmp/h0001.nc
// msrcp -period 365 ~/nco/data/in.nc mss:/ZENDER/tmp/h0002.nc
// msrcp -period 365 ~/nco/data/in.nc mss:/ZENDER/tmp/h0003.nc
// msrcp -period 365 ~/nco/data/in.nc mss:/ZENDER/tmp/h0004.nc

// WARNING: Changing values of variables below, especially coordinate variables, affects outcome of nco_tst.pl test script
// Other programs, e.g., ~/f/fff.F90, ~/c++/ccc.cc, ~/c/c.c may also break
// In particular, do not change number of elements in record coordinate, time, without simultaneously changing number of data in all record variables
// My (and NCO's) convention is that the _FillValue, if any, of any packed variable should be of the same type as the expanded variable. Hence _FillValue, add_offset, and scale_factor should all be of the same type. Variables that do not adhere to this convention are not supported.

// CDL Data constants:
// byte: 'a'
// char: "a"
// short: 1s
// int: 1 (no decimal point)
// float: 1.f (decimal point is required, f is required to distinguish from double)
// double: 1.0, 1.d, 1.0e-20 (decimal point is required, d is not required)
// 

// NCL usage:
// id_in=addfile("/home/zender/nco/data/in.nc","r")
// print(id_in)
// list_filevars(id_in)

netcdf in {
dimensions:
	dgn=1,bnd=2,lat=2,lat_grd=3,lev=3,rlev=3,lon=4,lon_grd=5,char_dmn_lng80=80,char_dmn_lng04=4,fl_dmn=3,lsmlev=6,wvl=2,time_udunits=3;lon_T42=128,lat_T42=64,lat_times_lon=8,gds_crd=8,lon_cal=10,lat_cal=10,time=unlimited;
variables:
	:Conventions = "CF-1.0";
	:history = "History global attribute.\n";
	:julian_day = 200000.04;
	:RCS_Header = "$Header: /data/zender/nco_20150216/nco/data/in.cdl,v 1.115 2010-08-09 18:11:55 zender Exp $";

	float lat(lat);
	lat:long_name = "Latitude (typically midpoints)";
	lat:units = "degrees_north";

	float lat_grd(lat_grd);
	lat_grd:long_name = "Latitude grid (typically interfaces)";
	lat_grd:units = "degrees_north";

	float lat_cpy(lat);
	float lev_cpy(lev);
	float lat_var(lat);
	float lat_wgt(lat);
	float lon_T42(lon_T42);
	float lat_T42(lat_T42);

	float lat_1D_rct(lat_times_lon);
	lat_1D_rct:long_name = "Latitude for 2D rectangular grid stored as 1D arrays";
	lat_1D_rct:units = "degrees_north";

	float lon_1D_rct(lat_times_lon);
	lon_1D_rct:long_name = "Longitude for 2D rectangular grid stored as 1D arrays";
	lon_1D_rct:units = "degrees_east";

	float lat_1D_rrg(lat_times_lon);
	lat_1D_rrg:long_name = "Latitude for 2D irregular grid stored as 1D arrays";
	lat_1D_rrg:units = "degrees_north";

	float lon_1D_rrg(lat_times_lon);
	lon_1D_rrg:long_name = "Longitude for 2D irregular grid stored as 1D arrays";
	lon_1D_rrg:units = "degrees_east";

	int lat_times_lon(lat_times_lon);
	lat_times_lon:long_name = "Element index (i.e., C-based storage order) for 2D coordinate grids stored as 1D arrays";

	float lat_2D_rct(lat,lon);
	lat_2D_rct:long_name = "Latitude for 2D rectangular grid stored as 2D array";
	lat_2D_rct:units = "degrees_north";

	float lon_2D_rct(lat,lon);
	lon_2D_rct:long_name = "Longitude for 2D rectangular grid stored as 2D array";
	lon_2D_rct:units = "degrees_east";

	float lat_2D_rrg(lat,lon);
	lat_2D_rrg:long_name = "Latitude for 2D irregular grid stored as 2D array";
	lat_2D_rrg:units = "degrees_north";

	float lon_2D_rrg(lat,lon);
	lon_2D_rrg:long_name = "Longitude for 2D irregular grid stored as 2D array";
	lon_2D_rrg:units = "degrees_east";

	int lat_times_lon_nbr;
	lat_times_lon_nbr:long_name = "Number of elements in 2D coordinate grids. Rectangular and irregular test grids have this many total elements. The coordinates and elements are stored as 1D or 2D arrays for grid types 1D and 2D respectively.";

	float lev(lev);
	lev:purpose = "Monotonically increasing coordinate pressure";
	lev:units = "hybrid_sigma_pressure";
	lev:positive = "down";
	lev:A_var = "hyam";
	lev:B_var = "hybm";
	lev:P0_var = "P0";
	lev:PS_var = "PS";
	lev:bounds = "ilev";

	float rlev(rlev);
	rlev:purpose = "Monotonically decreasing coordinate pressure";

	float lon(lon);
	lon:long_name = "Longitude (typically midpoints)";
	lon:units = "degrees_east";

	double lond(lon);
	lond:long_name = "Longitude (typically midpoints), double precision";
	lond:units = "degrees_east";

	float lonf(lon);
	lonf:long_name = "Longitude (typically midpoints), single precision";
	lonf:units = "degrees_east";

	float lon_grd(lon_grd);
	lon_grd:long_name = "Longitude grid (typically interfaces)";
	lon_grd:units = "degrees_east";

	double time(time);
	time: long_name = "time";
	time: units = "days since 1964-03-12 12:09:00 -9:00"; 
	time: calendar = "gregorian";


	double lon_cal(lon_cal);
	lon_cal: long_name = "lon_cal";
	lon_cal: units = "days since 1964-2-28"; 
	lon_cal: calendar = "365_day";


	double lat_cal(lat_cal);
	lat_cal: long_name = "lat_cal";
	lat_cal: units = "days since 1964-2-28"; 
	lat_cal: calendar = "360_day";


	float lsmlev(lsmlev);
	lsmlev:purpose = "Homebrew level coordinate for LSM";
	lsmlev:long_name = "Soil depth";
	lsmlev:units = "meter";
	float wvl(wvl);
	wvl:long_name = "Wavelength";
	wvl:units = "meter";

	int od(time);

	float area(lat);
	area:long_name = "area";
	area:units = "meter2";

	float hyam(lev);
	hyam:long_name = "hybrid A coefficient at layer midpoints";

	float hybm(lev);
	hybm:long_name = "hybrid B coefficient at layer midpoints";

	float P0;
	P0:long_name = "reference pressure";
	P0:units = "pascal";

	float cnv_CF_crd(gds_crd);
	cnv_CF_crd:long_name = "test CF coordinates conventions";
	cnv_CF_crd:coordinates = "lat_gds lon_gds ";
	cnv_CF_crd:reason = "Test whether coordinates attribute strings that end with a space break after nco_var_lst_crd_ass_add() call to nco_lst_prs_2d()";

	float PS(time,lat,lon);
	PS:long_name = "surface pressure";
	PS:units = "pascal";

	char fl_dmn(fl_dmn);
	fl_dmn:long_name = "Character coordinate";
	fl_dmn:units = "[chr]";

	double lat_gds(gds_crd);
	lat_gds:long_name = "Latitude";  
	lat_gds:standard_name = "latitude";
	lat_gds:units="degree";
	lat_gds:purpose = "1-D latitude coordinate referred to by geodesic grid variables";

	double lon_gds(gds_crd);
	lon_gds:long_name = "Longitude";
	lon_gds:standard_name = "longitude";
	lon_gds:units="degree";
	lon_gds:purpose = "1-D longitude coordinate referred to by geodesic grid variables";

	float gds_crd(gds_crd);
	gds_crd:long_name = "Geodesic coordinate";
	gds_crd:units = "degree";
	gds_crd:purpose = "enumerated coordinate like those that might define points in a geodesic grid";
	gds_crd:coordinates = "lat_gds lon_gds";

	float gds_var(gds_crd);
	gds_var:long_name = "Geodesic variable";
	gds_var:units = "meter";
	gds_var:purpose = "Test auxiliary coordinates like those that define geodesic grids";
	gds_var:coordinates = "lat_gds lon_gds";


	float gds_3dvar(time,gds_crd);
	gds_3dvar:long_name = "Geodesic variable";
	gds_3dvar:units = "meter";
	gds_3dvar:coordinates = "lat_gds lon_gds";
	gds_3dvar:purpose = "Test auxiliary coordinates like those that define geodesic grids";

	int nbdate;
	nbdate:long_name = "base date as 6- or 8-digit integer (YYMMDD or YYYYMMDD)";
	int date(time);
	date:long_name = "current date as 6- or 8-digit integer (YYMMDD or YYYYMMDD)";

	float lon_wgt(lon);
	lon_wgt:long_name = "Gaussian weights";
	lon_wgt:purpose = "Gaussian weights which sum to two for n = 4. These weights are all have floor of 0.0 so should cause SIGFPE when applied to integer types in weighted average.";

	float msk_prt_mss_prt(lon);
	msk_prt_mss_prt:long_name = "partial mask, partial missing value example";
	msk_prt_mss_prt:_FillValue = 1.0e36f;

	float mss_val(lon);
	mss_val:long_name = "partial missing value example";
	mss_val:_FillValue = 1.0e36f;

	float mss_val_scl;
	mss_val_scl:long_name = "scalar missing value";
	mss_val_scl:_FillValue = 1.0e36f;

	float mss_val_fst(lon);
	mss_val_fst:long_name = "offset partial missing value example";
	mss_val_fst:_FillValue = -999.0f;

	float fll_val(lon);
	fll_val:long_name = "_FillValue example";
	fll_val:_FillValue = -999.0f;

	float fll_val_mss_val(lon);
	fll_val_mss_val:long_name = "_FillValue example";
	fll_val_mss_val:_FillValue = -999.0f;
	fll_val_mss_val:missing_value = -999.0f;

	float nm_spc;
	nm_spc:long_name = "Variable name with space (invalid)";

	float nm_pnd;
	nm_pnd:long_name = "Variable name with pound symbol (invalid)";

	float no_mss_val(lon);
	no_mss_val:long_name = "no missing value";

	float val_one_mss(lat);
	val_one_mss:long_name = "one regular value, one missing value";
	val_one_mss:_FillValue = 1.0e36f;

	short pck;
	pck:long_name = "Packed scalar variable";
	pck:note = "Original packed value was 1s with scale_factor = 2.0d and add_offset = 1.0d. Unpacked value should be 3.0 = 2.0d*1s + 1.0d. NCO algorithms would pack this variable as scale_factor = 0.0d and add_offset = 3.0d.";
	pck:scale_factor = 2.0d;
	pck:add_offset = 1.0d;

	short pck_arr(lon);
	pck_arr:long_name = "Packed array";
	pck_arr:note = "Packed value is -32767s, 0s, 1s, 32767s, unpacked is same in double";
	pck_arr:scale_factor = 1.0d;
	pck_arr:add_offset = 0.0d;

	double upk;
	upk:long_name = "Unpacked scalar variable";
	upk:note = "Unpacked value is 3.0d0, upk=unpack(pck)= 2.0d0*1s + 1.0d0 = 3.0d0. Packing this variable should create an NC_SHORT scalar = 0s with packing attribute add_offset=3.0d and either no scale_factor (ncap) or scale_factor = 0.0d (ncpdq).";

	double upk_arr(lon);
	upk_arr:long_name = "Unpacked array";
	upk_arr:note = "Unpacked value is -32767.d, 0.d, 1.d, 32767.d, packed is same in short. Packing algorithm should yield an NC_SHORT array = [] with packing attributes scale_factor=1.0d, add_offset=0.0d";

	int val_one_int;
	val_one_int:long_name = "scalar equal to 1";
	val_one_int:_FillValue = -99l;

	int val_one_one_int(lat);
	val_one_one_int:long_name = "1, 1";
	val_one_one_int:_FillValue = -99l;

	short val_max_max_sht(lat);
	val_max_max_sht:long_name = "17000, 17000";
	val_max_max_sht:_FillValue = -99s;

	int val_one_mss_int(lat);
	val_one_mss_int:long_name = "1, mss_val";
	val_one_mss_int:_FillValue = -99l;

	float val_half;
	val_half:long_name = "Scalar with value 0.5";
	val_half:_FillValue = 1.0e36f;

	float val_half_half(lat);
	val_half_half:long_name = "0.5,0.5";
	val_half_half:_FillValue = 1.0e36f;

	float wgt_one(lat);
	wgt_one:long_name = "all values are one";

	float mss_val_all(lon);
	mss_val_all:long_name = "all missing values example";
	mss_val_all:_FillValue = 1.0e36f;

	float scalar_var;
	scalar_var:long_name = "scalar variable";
	scalar_var:units = "fraction";

	float float_var;
	float_var:long_name = "float";

	double double_var;
	double_var:long_name = "double";

	double double_var2;
	double_var2:long_name = "double";
	double_var2:_FillValue = 1.0e36;

	double pi;
	pi:long_name = "Pi";
	pi:units = "fraction";

	int int_var;
	int_var:long_name = "int";

	short short_var;
	short_var:long_name = "short";

	char char_var;
	char_var:long_name = "char";

	char char_var_space;
	char_var_space:long_name = "Character variable with whitespace on ends";

	char char_var_nul;
	char_var_nul:long_name = "Character variable containing one NUL";

	char char_var_multinul(lev);
	char_var_multinul:long_name = "Character variable containing multiple NULs";

	char fl_nm(char_dmn_lng80);
	fl_nm:long_name = "Variable contains a file name";

	char fl_nm_arr(fl_dmn,char_dmn_lng80);
	fl_nm_arr:long_name = "Variable that contains a short array of file names";
	fl_nm_arr:units = "[sng]";

	char non_nul_trm_char_one_dmn(char_dmn_lng04);
	non_nul_trm_char_one_dmn:long_name = "Variable contains a one-dimensional array of characters that is not NUL-terminated";
	non_nul_trm_char_one_dmn:units = "[chr]";

	char non_nul_trm_char_two_dmn(fl_dmn,char_dmn_lng04);
	non_nul_trm_char_two_dmn:long_name = "Variable contains a two-dimensional array of characters that are not NUL-terminated";
	non_nul_trm_char_two_dmn:units = "[chr]";

	byte byte_var;
	byte_var:long_name = "byte";

	byte byte_var_neg;
	byte_var_neg:long_name = "negative byte";

	float zero;
	zero:long_name = "zero";

	float one;
	one:long_name = "one";

	float two;
	two:long_name = "two";

	double e_dbl;
	e_dbl:long_name = "e, natural logarithm base";

	float e_flt;
	e_flt:long_name = "e, natural logarithm base";

	float three;
	three:long_name = "three";

	float four;
	four:long_name = "four";

	float negative_one;
	negative_one:long_name = "negative one";

	float lev_var(lev);
	lev_var:long_name = "lev_var";

	float lev_wgt(lev);
	lev_wgt:long_name = "lev_wgt";

	float g;
	g:long_name = "g";

	float z(lev);
	z:long_name = "Height";
	z:units = "meter";
	z:purpose = "Height stored with a monotonically increasing coordinate";

	float rz(rlev);
	rz:long_name = "Height";
	rz:units = "meter";
	rz:purpose = "Height stored with a monotonically decreasing coordinate";

	float one_dmn_var(bnd);

	int one_dmn_int_val_one(lat);
	int one_dmn_int_val_two(lat);

	float att_var;
	att_var:byte_att = '\0';
	att_var:char_att = "Sentence one.\nSentence two.\n";
	att_var:short_att = 37s;
	att_var:int_att = 73l;
	att_var:float_att = 73.0f,72.0f,71.0f;
	att_var:double_att = 73.0d;

	int bnd_var(lev,bnd);
	bnd_var:byte_att = '\0';
	bnd_var:char_att = "Sentence one.\nSentence two.\n";
	bnd_var:short_att = 37s;
	bnd_var:int_att = 73;
	bnd_var:float_att = 73.f;
	bnd_var:double_att = 73.d;

	float three_dmn_var(lat,lev,lon);
	three_dmn_var:long_name = "three dimensional variable with CCM coordinate convention C=[lat,lev,lon], Fortran=(lon,lev,lat)";
	three_dmn_var:units = "fraction";

	float three_dmn_var_crd(lev,lat,lon);
	three_dmn_var_crd:long_name = "three dimensional variable with COORDS coordinate convention C=[lev,lat,lon], Fortran=(lon,lat,lev)";
	three_dmn_var_crd:units = "fraction";

	float prs_sfc(time,lat,lon);
	prs_sfc:long_name = "Surface pressure";
	prs_sfc:units = "pascal";

	float H2O;
	float H2OH2O;
	float H2SO4;
	float H2O_lqd;
	float H2O_ice;
	float Q;
	float Q1;
	float AQ01;
	float QQ01;
	float QA01;
	float Q01Q;
	float Q01;
	float Q02;
	float Q03;
	float Q04;
	float Q05;
	float Q06;
	float Q07;
	float Q08;
	float Q09;
	float Q10;
	float Q11;
	float Q12;
	float Q13;
	float Q14;
	float Q15;
	float Q16;
	float Q17;
	float Q18;
	float Q19;
	float Q20;
	float Q21;
	float Q22;
	float Q23;
	float Q24;
	float Q25;
	float Q26;
	float Q27;
	float Q28;
	float Q29;
	float Q30;
	float Q31;
	float Q32;
	float Q33;
	float Q34;
	float Q35;
	float Q36;
	float Q37;
	float Q38;
	float Q39;
	float Q40;
	float Q41;
	float Q42;
	float Q43;
	float Q44;
	float Q45;
	float Q46;
	float Q47;
	float Q48;
	float Q49;
	float Q50;
	float Q51;
	float Q52;
	float Q53;
	float Q54;
	float Q55;
	float Q56;
	float Q57;
	float Q58;
	float Q59;
	float Q60;
	float Q61;
	float Q62;
	float Q63;
	float Q64;
	float Q65;
	float Q66;
	float Q67;
	float Q68;
	float Q69;
	float Q70;
	float Q71;
	float Q72;
	float Q73;
	float Q74;
	float Q75;
	float Q76;
	float Q77;
	float Q78;
	float Q79;
	float Q80;
	float Q81;
	float Q82;
	float Q83;
	float Q84;
	float Q85;
	float Q86;
	float Q87;
	float Q88;
	float Q89;
	float Q90;
	float Q91;
	float Q92;
	float Q93;
	float Q94;
	float Q95;
	float Q96;
	float Q97;
	float Q98;
	float Q99;
	float Q100;

	float two_dmn_var(lat,lev);
	two_dmn_var:long_name = "two dimensional variable";
	two_dmn_var:units = "fraction";

	float var_msk(lat,lon);
	var_msk:long_name = "Float field for testing masks and wheres";
	var_msk:units = "fraction";

	float mask(lat,lon);
	mask:long_name = "Purpose is to mask a variable like ORO";
	mask:units = "fraction";

	float ORO(lat,lon);
	ORO:long_name = "Orography, an enumerated yet continuous type: ocean=0.0, land=1.0, sea ice=2.0";
	ORO:units = "fraction";

	float weight(lat);
	weight:long_name = "Gaussian weight";
	weight:units = "fraction";

	float gw(lat);
	gw:long_name = "gw variable like gw";
	gw:units = "fraction";

	float gw_T42(lat_T42);
	gw_T42:long_name = "gw variable like gw_T42";
	gw_T42:units = "fraction";

	float rec_var_flt(time);
	rec_var_flt:long_name = "record variable, float";

	double rec_var_dbl(time);
	rec_var_dbl:long_name = "record variable, double";

	int one_dmn_rec_var(time);
	one_dmn_rec_var:long_name = "one dimensional record variable";
	one_dmn_rec_var:units = "second";
        
	int RDM(time);
        
	float tpt(time);
	tpt:long_name = "Temperature";
	tpt:units = "kelvin";
	tpt:hieght = "Leave hieght mispelled for NCO User's guide example";

	double rec_var_dbl_mss_val_dbl_upk(time);
	rec_var_dbl_mss_val_dbl_upk:long_name = "record variable, double, with double missing values";
	rec_var_dbl_mss_val_dbl_upk:purpose = "This variable is used to generate the packed variable rec_var_dbl_mss_val_dbl_pck, so its _FillValue should not be too far out of range, i.e., it should be representable by a short. However, the _FillValue should itself be the same type as the unpacked variable, NC_DOUBLE in this case.";
	rec_var_dbl_mss_val_dbl_upk:_FillValue = -999.;

	short rec_var_dbl_mss_val_dbl_pck(time);
	rec_var_dbl_mss_val_dbl_pck:long_name = "record variable, double, with double missing values, packed";
	rec_var_dbl_mss_val_dbl_pck:purpose = "Packed version of rec_var_dbl_mss_val_dbl_upk";
	rec_var_dbl_mss_val_dbl_pck:_FillValue = -999s;
	rec_var_dbl_mss_val_dbl_pck:missing_value = -999.;
        rec_var_dbl_mss_val_dbl_pck:scale_factor = -9.15541313801785e-05;
        rec_var_dbl_mss_val_dbl_pck:add_offset = 5. ;

	short scl_dbl_pck;
	scl_dbl_pck:long_name = "scalar variable, double, packed";
	scl_dbl_pck:purpose = "Packed version of number with ncdiff subtraction bug";
        scl_dbl_pck:scale_factor = -9.15541313801785e-05;
        scl_dbl_pck:add_offset = 5. ;

	float rec_var_flt_mss_val_flt(time);
	rec_var_flt_mss_val_flt:long_name = "record variable, float, with float missing values";
	rec_var_flt_mss_val_flt:_FillValue = 1.0e36f;

	float rec_var_flt_mss_val_flt_all(time);
	rec_var_flt_mss_val_flt_all:long_name = "record variable, float, with float missing values in every position";
	rec_var_flt_mss_val_flt_all:_FillValue = 1.0e36f;

	float rec_var_flt_mss_val_flt_all_but_one(time);
	rec_var_flt_mss_val_flt_all_but_one:long_name = "record variable, float, with float missing values in every position but one";
	rec_var_flt_mss_val_flt_all_but_one:_FillValue = 1.0e36f;

	float rec_var_flt_mss_val_flt_all_but_two(time);
	rec_var_flt_mss_val_flt_all_but_two:long_name = "record variable, float, with float missing values in every position but two";
	rec_var_flt_mss_val_flt_all_but_two:_FillValue = 1.0e36f;

	short rec_var_flt_pck(time);
	rec_var_flt_pck:long_name = "record variable, float, packed";
        rec_var_flt_pck:purpose = "Demonstrate that rounding of means of packed data are handled correctly";
        rec_var_flt_pck:scale_factor = 0.1f;
        rec_var_flt_pck:add_offset = 100.0f;

	short rec_var_dbl_pck(time);
	rec_var_dbl_pck:long_name = "record variable, double, packed";
        rec_var_dbl_pck:purpose = "Demonstrate that rounding of means of packed data are handled correctly";
        rec_var_dbl_pck:scale_factor = 0.1;
		rec_var_dbl_pck:add_offset = 100.0;
	
	short non_rec_var_flt_pck(lon);
		non_rec_var_flt_pck:long_name = "regular variable, float, packed";
        non_rec_var_flt_pck:purpose = "Demonstrate that non-rec dim packed vars are handled correctly";
        non_rec_var_flt_pck:scale_factor = 0.1f;
        non_rec_var_flt_pck:add_offset = 100.0f;

	float rec_var_flt_mss_val_dbl(time);
	rec_var_flt_mss_val_dbl:long_name = "record variable, float, with double missing values";
	rec_var_flt_mss_val_dbl:_FillValue = 1.0e36f;
	rec_var_flt_mss_val_dbl:missing_value = 1.0e36;
	rec_var_flt_mss_val_dbl:note = "The correct average of this variable is 5.0";

	float rec_var_flt_mss_val_int(time);
	rec_var_flt_mss_val_int:long_name = "record variable, float, with integer missing values";
	rec_var_flt_mss_val_int:_FillValue = -999.0f;
	rec_var_flt_mss_val_int:missing_value = -999;

	int rec_var_int_mss_val_int(time);
	rec_var_int_mss_val_int:long_name = "record variable, integer, with integer missing values";
	rec_var_int_mss_val_int:_FillValue = -999;

	int rec_var_int_mss_val_flt(time);
	rec_var_int_mss_val_flt:long_name = "record variable, integer, with float missing values";
	rec_var_int_mss_val_flt:_FillValue = -999;
	rec_var_int_mss_val_flt:missing_value = -999.0f;

	int rec_var_int_mss_val_dbl(time);
	rec_var_int_mss_val_dbl:long_name = "record variable, integer, with double missing values";
	rec_var_int_mss_val_dbl:_FillValue = -999;
	rec_var_int_mss_val_dbl:missing_value = -999.0;

	int rec_var_dbl_mss_val_dbl_pck_lng(time);
	rec_var_dbl_mss_val_dbl_pck_lng:long_name = "record variable, double packed as long, with double missing values";
	rec_var_dbl_mss_val_dbl_pck_lng:purpose = "although not usual, packing doubles into longs (rather than shorts) is still a considerable cost savings";
	rec_var_dbl_mss_val_dbl_pck_lng:_FillValue = -999;
	rec_var_dbl_mss_val_dbl_pck_lng:missing_value = -999.0;
        rec_var_dbl_mss_val_dbl_pck_lng:scale_factor = -9.15541313801785e-05 ;
        rec_var_dbl_mss_val_dbl_pck_lng:add_offset = 5. ;

	char one_dmn_rec_var_sng(time);
	one_dmn_rec_var_sng:long_name = "one dimensional record variable of string";

	float time_lon(time,lon);
	time_lon:long_name = "Record variable of longitude coordinate";

	char two_dmn_rec_var_sng(time,lev);
	two_dmn_rec_var_sng:long_name = "two dimensional record variable of string";

	float two_dmn_rec_var(time,lev);
	two_dmn_rec_var:long_name = "two dimensional record variable";
	two_dmn_rec_var:units = "watt meter-2";

	float three_dmn_rec_var(time,lat,lon);
	three_dmn_rec_var:long_name = "three dimensional record variable";
	three_dmn_rec_var:units = "watt meter-2";

	double three_dmn_var_dbl(time,lat,lon);
	three_dmn_var_dbl:long_name = "three dimensional record variable of type double";
	three_dmn_var_dbl:units = "watt meter-2";
	three_dmn_var_dbl:_FillValue = -99. ;

	int three_dmn_var_int(time,lat,lon);
	three_dmn_var_int:long_name = "three dimensional record variable of type int";
	three_dmn_var_int:units = "watt meter-2";
	three_dmn_var_int:_FillValue = -99 ;
	
	short three_dmn_var_sht(time,lat,lon);
	three_dmn_var_sht:long_name = "three dimensional record variable";
	three_dmn_var_sht:units = "watt meter-2";
	three_dmn_var_sht:_FillValue = -99s ;


	int th(time,lat,lon);
	th:long_name = "three dimensional record variable";
	th:units = "watt meter-2";
	th:_FillValue = -99;


	float td(time,dgn);
	td:long_name = "two dimensional record variable stored in td (time,dgn) order (dgn means degenerate, i.e., of size 1)";

	float tx(time,lon);
	tx:long_name = "two dimensional record variable stored in tx (time,lon) order";

	float ty(time,lat);
	ty:long_name = "two dimensional record variable stored in ty (time,lat) order";

	float tz(time,lev);
	tz:long_name = "two dimensional record variable stored in tz (time,lev) order";

	float txyz(time,lon,lat,lev);
	txyz:long_name = "four dimensional record variable stored in txyz (time,lon,lat,lev) order";


	float four_dmn_rec_var(time,lat,lev,lon);
	four_dmn_rec_var:long_name = "four dimensional record variable";
	four_dmn_rec_var:units = "watt meter-2";

//	double three_double_dmn(time,lon,lon);
	
	double time_udunits(time_udunits);
	time_udunits:units = "hours since 1900-01-01 00:00:0.0";
	time_udunits:delta_t = "0000-00-00 06:00:0.0";

	float u(time);
	u:long_name = "Zonal wind speed";
	u:units = "meter second-1";

	float v(time);
	v:long_name = "Meridional wind speed";
	v:units = "meter second-1";

	float var_1D_rct(lat_times_lon);
	var_1D_rct:long_name = "Variable for 2D rectangular grid stored as 1D arrays";

	float var_1D_rrg(lat_times_lon);
	var_1D_rrg:long_name = "Variable for 2D irregular grid stored as 1D arrays";

	float var_2D_rct(lat,lon);
	var_2D_rct:long_name = "Variable for 2D rectangular grid stored as 2D array";

	float var_2D_rrg(lat,lon);
	var_2D_rrg:long_name = "Variable for 2D irregular grid stored as 2D array";

	float var_nm-dash;
	var_nm-dash:long_name = "Variable and attribute names include dash characters";
	var_nm-dash:att_nm-dash = 1.0e36f;

	float var_nm.dot;
	var_nm.dot:long_name = "Variable and attribute names include dot characters";
//	20070102: Periods in attribute names choke OPeNDAP from FC7 RPM TODO nco911
//	20091105: Periods in attribute names choke ncgen   from RHEL5   TODO nco911
//	var_nm.dot:att_nm.dot = 1.0e36f;

	float wnd_spd(time,lat,lon);
	wnd_spd:long_name = "wind speed";
	wnd_spd:units = "meter second-1";
	wnd_spd:_FillValue = -999.0f;

data:
	att_var=10.;
	area=10.,10.;
	bnd_var=1,2,3,4,5,6;
	byte_var='z';
	byte_var_neg=-122;
	char_var="z";
	char_var_multinul="\b\n\0";
	char_var_nul='\0';
	char_var_space=" ";
	cnv_CF_crd=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8;
	double_var=10.;
	double_var2=10.;
	e_dbl=2.71828182846;
	e_flt=2.71828182846;
// 	20100809: Single quotes around NC_CHAR coordinates required as of 4.1.2-beta1-snapshot2010080820
// 	20100809: Double quotes cause "String constant too long" error in ncgen
	fl_dmn='a','b','3';
	fl_nm="/home/zender/nco/data/in.cdl";
	float_var=10.;
	four=4.;
	g=9.8;
	gw=10.,10.;
	gw_T42=-87.863799,-85.096527,-82.312913,-79.525607,-76.736900,-73.947515,-71.157752,-68.367756,-65.577607,-62.787352,-59.997020,-57.206632,-54.416200,-51.625734,-48.835241,-46.044727,-43.254195,-40.463648,-37.673090,-34.882521,-32.091944,-29.301360,-26.510769,-23.720174,-20.929574,-18.138971,-15.348365,-12.557756,-9.767146,-6.976534,-4.185921,-1.395307,1.395307,4.185921,6.976534,9.767146,12.557756,15.348365,18.138971,20.929574,23.720174,26.510769,29.301360,32.091944,34.882521,37.673090,40.463648,43.254195,46.044727,48.835241,51.625734,54.416200,57.206632,59.997020,62.787352,65.577607,68.367756,71.157752,73.947515,76.736900,79.525607,82.312913,85.096527,87.863799;
	hyam=0.0802583,0.0438226,0.0;
	hybm=0.0187849,0.457453,0.992528;
	P0=100000;
	gds_crd=0,1,2,3,4,5,6,7;
	gds_var=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8;
	gds_3dvar=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8,
	          274.1,274.2,274.3,274.4,274.5,274.6,274.7,274.8,
	          275.1,275.2,275.3,275.4,275.5,274.5,275.7,275.8,
	          276.1,276.2,276.3,276.4,276.5,276.5,276.7,276.8,
	          277.1,277.2,277.3,277.4,277.5,277.5,277.7,277.8,
	          278.1,278.2,278.3,278.4,278.5,278.6,278.7,278.8,
	          279.1,279.2,279.3,279.4,279.5,279.9,279.7,279.8,
	          280.1,280.2,280.3,280.4,280.5,280.9,280.7,280.8,
	          281.1,281.2,281.3,281.4,281.5,281.9,281.7,281.8,
	          282.1,282.2,282.3,282.4,282.5,282.9,282.7,282.8;
	lat_gds=-90, -30,  -30,    0,   0, 30,  30,  90;
	lon_gds=  0,   0,  180,    0, 180,  0, 180,   0;
	lat=-90,90;
        lat_cal=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	lon_cal=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	lat_times_lon=0,1,2,3,4,5,6,7;
	lat_times_lon_nbr=8;
	lat_1D_rct=-90, -90,  -90,  -90,  90, 90,  90,  90;
	lon_1D_rct=  0,  90,  180,  270,   0, 90, 180, 270;
	lat_1D_rrg=-90, -30,  -30,    0,   0, 30,  30,  90;
	lon_1D_rrg=  0,   0,  180,    0, 180,  0, 180,   0;
	lat_2D_rct=-90, -90,  -90,  -90,  90, 90,  90,  90;
	lon_2D_rct=  0,  90,  180,  270,   0, 90, 180, 270;
	lat_2D_rrg=-90, -30,  -30,    0,   0, 30,  30,  90;
	lon_2D_rrg=  0,   0,  180,    0, 180,  0, 180,   0;
	lat_grd=-90,0,90;
	lat_cpy=-90,90;
	lat_var=1.,2.;
	lat_wgt=1.,2.;
//	lat_T42=0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63;
	lat_T42=-88.240089,-85.092445,-82.311981,-79.525253,-76.736732,-73.947418,-71.157700,-68.367722,-65.577576,-62.787331,-59.997005,-57.206619,-54.416191,-51.625729,-48.835236,-46.044724,-43.254192,-40.463646,-37.673088,-34.882519,-32.091942,-29.301357,-26.510769,-23.720173,-20.929573,-18.138969,-15.348364,-12.557755,-9.767145,-6.976533,-4.185921,-1.395307,1.395307,4.185921,6.976533,9.767145,12.557755,15.348364,18.138969,20.929573,23.720173,26.510769,29.301357,32.091942,34.882519,37.673088,40.463646,43.254192,46.044724,48.835236,51.625729,54.416191,57.206619,59.997005,62.787331,65.577576,68.367722,71.157700,73.947418,76.736732,79.525253,82.311981,85.092445,88.240089;
	lsmlev=0.05,0.1,0.2,0.5,1.0,3.0;
	lev=100,500,1000;
	lev_cpy=100,500,1000;
	lev_var=100.,500.,1000.;
	lev_wgt=10,2,1;
	lon=0,90,180,270;
	lond=0,90,180,270;
	lonf=0,90,180,270;
	lon_grd=-45,45,135,225,315;
	lon_wgt=0.347855,0.652145,0.652145,0.347855;
//	lon_T42=0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127;
	lon_T42=0.000000,2.812500,5.625000,8.437500,11.250000,14.062500,16.875000,19.687500,22.500000,25.312500,28.125000,30.937500,33.750000,36.562500,39.375000,42.187500,45.000000,47.812500,50.625000,53.437500,56.250000,59.062500,61.875000,64.687500,67.500000,70.312500,73.125000,75.937500,78.750000,81.562500,84.375000,87.187500,90.000000,92.812500,95.625000,98.437500,101.250000,104.062500,106.875000,109.687500,112.500000,115.312500,118.125000,120.937500,123.750000,126.562500,129.375000,132.187500,135.000000,137.812500,140.625000,143.437500,146.250000,149.062500,151.875000,154.687500,157.500000,160.312500,163.125000,165.937500,168.750000,171.562500,174.375000,177.187500,180.000000,182.812500,185.625000,188.437500,191.250000,194.062500,196.875000,199.687500,202.500000,205.312500,208.125000,210.937500,213.750000,216.562500,219.375000,222.187500,225.000000,227.812500,230.625000,233.437500,236.250000,239.062500,241.875000,244.687500,247.500000,250.312500,253.125000,255.937500,258.750000,261.562500,264.375000,267.187500,270.000000,272.812500,275.625000,278.437500,281.250000,284.062500,286.875000,289.687500,292.500000,295.312500,298.125000,300.937500,303.750000,306.562500,309.375000,312.187500,315.000000,317.812500,320.625000,323.437500,326.250000,329.062500,331.875000,334.687500,337.500000,340.312500,343.125000,345.937500,348.750000,351.562500,354.375000,357.187500;
	mask=0.,1.,0.,0.,1.,1.,0.,2.;
	var_msk=0.,1.,0.,0.,1.,1.,0.,2.;
	ORO=0.,1.,0.,0.,1.,1.,0.,2.;
//	mask=0.,0.,0.,0.,0.,0.,0.,0.;
//	mask=1.,1.,1.,1.,1.,1.,1.,1.;
	fll_val=73,-999,73,-999;
	fll_val_mss_val=73,-999,73,-999;
	msk_prt_mss_prt=0.5,1.0e36,1.5,1.0e36;
	mss_val=73,1.0e36,73,1.0e36;
	mss_val_all=1.0e36,1.0e36,1.0e36,1.0e36;
	mss_val_fst=-999,73,-999,73;
	mss_val_scl=1.0e36;
	negative_one=-1.;
	nm_pnd=1;
	nm_spc=1;
	no_mss_val=73,1.0e36,73,1.0e36;
	non_nul_trm_char_one_dmn='a','b';
	non_nul_trm_char_two_dmn="abcd","efgh","ijkm";
	one=1.;
	one_dmn_rec_var=1,2,3,4,5,6,7,8,9,10;
	RDM=1,9,36,84,126,126,84,36,9,1;
	one_dmn_rec_var_sng="Hello Wor";
	one_dmn_var=1.,10.;
	one_dmn_int_val_one=1,1;
	one_dmn_int_val_two=2,2;
	pck=1;
	pck_arr=-32767,0,1,32767;
	pi=3.1415926535897932384626433832795029;
	upk=3.;
	upk_arr=-32767.,0.,1.,32767.;
	H2O=1.0;
	H2OH2O=1.0;
	H2SO4=1.0;
	H2O_lqd=1.0;
	H2O_ice=1.0;
	Q=1.0e36;
	Q1=1.0e36;
	AQ01=1.0e36;
	QQ01=1.0e36;
	QA01=1.0e36;
	Q01Q=1.0e36;
	Q01=1;
	Q02=2;
	Q03=3;
	Q04=4;
	Q05=5;
	Q06=6;
	Q07=7;
	Q08=8;
	Q09=9;
	Q10=10;
	Q11=11;
	Q12=12;
	Q13=13;
	Q14=14;
	Q15=15;
	Q16=16;
	Q17=17;
	Q18=18;
	Q19=19;
	Q20=20;
	Q21=21;
	Q22=22;
	Q23=23;
	Q24=24;
	Q25=25;
	Q26=26;
	Q27=27;
	Q28=28;
	Q29=29;
	Q30=30;
	Q31=31;
	Q32=32;
	Q33=33;
	Q34=34;
	Q35=35;
	Q36=36;
	Q37=37;
	Q38=38;
	Q39=39;
	Q40=40;
	Q41=41;
	Q42=42;
	Q43=43;
	Q44=44;
	Q45=45;
	Q46=46;
	Q47=47;
	Q48=48;
	Q49=49;
	Q50=50;
	Q51=51;
	Q52=52;
	Q53=53;
	Q54=54;
	Q55=55;
	Q56=56;
	Q57=57;
	Q58=58;
	Q59=59;
	Q60=60;
	Q61=61;
	Q62=62;
	Q63=63;
	Q64=64;
	Q65=65;
	Q66=66;
	Q67=67;
	Q68=68;
	Q69=69;
	Q70=70;
	Q71=71;
	Q72=72;
	Q73=73;
	Q74=74;
	Q75=75;
	Q76=76;
	Q77=77;
	Q78=78;
	Q79=79;
	Q80=80;
	Q81=81;
	Q82=82;
	Q83=83;
	Q84=84;
	Q85=85;
	Q86=86;
	Q87=87;
	Q88=88;
	Q89=89;
	Q90=90;
	Q91=91;
	Q92=92;
	Q93=93;
	Q94=94;
	Q95=95;
	Q96=96;
	Q97=97;
	Q98=98;
	Q99=99;
	Q100=100;
	rec_var_dbl=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	rec_var_flt=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	rec_var_flt_pck=1,2,3,4,5,6,7,8,9,10;
	rec_var_dbl_pck=1,2,3,4,5,6,7,8,9,10;
	non_rec_var_flt_pck=1,2,3,4;
	rec_var_dbl_mss_val_dbl_pck=-999,32767,21845,10922,0,-10922,-21845,-32767,-999,-999;
	rec_var_dbl_mss_val_dbl_upk=-999.,2.,3.,4.,5.,6.,7.,8.,-999.,-999.;
	rec_var_flt_mss_val_dbl=1.0e36,2.,3.,4.,5.,6.,7.,8.,1.0e36,1.0e36;
	rec_var_flt_mss_val_flt=1.0e36,2.,3.,4.,5.,6.,7.,8.,1.0e36,1.0e36;
	rec_var_flt_mss_val_flt_all=1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36;
	rec_var_flt_mss_val_flt_all_but_one=1.0e36,1.0e36,1.0e36,1.0e36,5.0,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36;
	rec_var_flt_mss_val_flt_all_but_two=1.0e36,1.0e36,1.0e36,1.0e36,5.0,1.0e36,1.0e36,1.0e36,1.0e36,10.0;
	rec_var_flt_mss_val_int=-999.,2.,3.,4.,5.,6.,7.,8.,-999.,-999.;
	rec_var_int_mss_val_int=-999,2,3,4,5,6,7,8,-999,-999;
	rec_var_int_mss_val_flt=-999,2,3,4,5,6,7,8,-999,-999;
	rec_var_dbl_mss_val_dbl_pck_lng=-999,32767,21845,10922,0,-10922,-21845,-32767,-999,-999;
	rec_var_int_mss_val_dbl=-999,2,3,4,5,6,7,8,-999,-999;
	rlev=1000,500,100;
	rz=0,5000,17000;
	scl_dbl_pck=10922;
	scalar_var=10.;
	short_var=10;
	three=3.;
	three_dmn_var=0.,1.,2.,3.,4.,5.,6.,7.,8.,9.,10.,11.,12.,13.,14.,15.,16.,17.,18.,19.,20.,21.,22.,23.;
	three_dmn_var_crd=0.,1.,2.,3.,12.,13.,14.,15.,4.,5.,6.,7.,16.,17.,18.,19.,8.,9.,10.,11.,20.,21.,22.,23.;
	time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	od=20,22,24,26,28,30,32,34,36,38 ;
	tpt=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8,273.9,274.0;
	two=2.;
	two_dmn_var=1.5,5.5,9.5,13.5,17.5,21.5;
	u=1.,0.,1.,0.,1.,0.,1.,0.,1.,0.;
	v=0.,1.,0.,1.,0.,1.,0.,1.,0.,1.;
	val_half=0.5;
	val_half_half=0.5,0.5;
	val_max_max_sht=17000,17000;
	val_one_int=1;
	val_one_mss=1.,1.0e36;
	val_one_mss_int=1,-99;
	val_one_one_int=1,1;
	var_nm-dash=1.0;
	var_nm.dot=1.0;
	var_1D_rct=0.,1.,0.,0.,1.,1.,0.,2.;
	var_1D_rrg=0.,1.,0.,0.,1.,1.,0.,2.;
	var_2D_rct=0.,1.,0.,0.,1.,1.,0.,2.;
	var_2D_rrg=0.,1.,0.,0.,1.,1.,0.,2.;
	weight=10.,10.;
	wgt_one=1.,1.;
	wvl=0.5e-6,1.0e-6;
	z=17000,5000,0;
	zero=0.;
 	date=640312,640313,640314,640315,640316,640317,640318,640319,640320,640321;
 	int_var=10;
 	nbdate=640312;
	fl_nm_arr="/data/zender/dstccm04/dstccm04_8589_01.nc",
		"/data/zender/dstccm04/dstccm04_8589_02.nc",
		"/data/zender/dstccm04/dstccm04_8589_03.nc";
	time_lon=0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0;
	two_dmn_rec_var_sng="abc",
				"bcd",
				"cde",
				"def",
				"efg",
				"fgh",
				"ghi",
				"hij",
				"jkl",
				"klm";
	two_dmn_rec_var=1.,2.0,3.,
			1.,2.1,3.,
			1.,2.2,3.,
			1.,2.3,3.,
			1.,2.4,3.,
			1.,2.5,3.,
			1.,2.6,3.,
			1.,2.7,3.,
			1.,2.8,3.,
			1.,2.9,3.;
	three_dmn_rec_var= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
  				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				73,74,75,76,77,78,79,80;
	prs_sfc=		 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
  				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				73,74,75,76,77,78,79,80;
	PS=			101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
  				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325;
	three_dmn_var_dbl= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				-99,-99,-99,-99,-99,-99,-99,-99,
				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				-99,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				-99,74,75,76,77,78,79,-99;
	three_dmn_var_int= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				-99,-99,-99,-99,-99,-99,-99,-99,
				25,26,27,28,29,30,31,32,
				33,34,35,36,37,38,39,40,
				41,-99,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				-99,58,59,60,-99,62,63,64,
				65,-99,67,68,69,70,71,72,
				-99,74,75,-99,77,78,79,80;
	three_dmn_var_sht= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 -99,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
				-99,34,35,-99,37,38,39,40,
				41,42,43,44,-99,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,-99,61,62,63,64,
				65,66,67,68,69,70,71,72,
				-99,-99,-99,-99,-99,-99,-99,-99;
	th=			1, 2, 3, 4, 5, 6, 7, 8,
				9,10,11,12,13,14,15,16,
			  	17,18,19,20,21,22,23,24,
			  	-99,-99,-99,-99,-99,-99,-99,-99,
			  	33,34,35,36,37,38,39,40,
			  	41,42,43,44,45,46,47,48,
			  	49,50,51,52,53,54,55,56,
			  	-99,58,59,60,61,62,63,64,
			  	65,66,67,68,69,70,71,72,
			 	-99,74,75,76,77,78,79,-99;
	four_dmn_rec_var= 	  1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12,
				 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24,
				 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36,
				 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48,
				 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60,
				 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72,
				 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84,
				 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96,
				 97, 98, 99,100,101,102,103,104,105,106,107,108,
				109,110,111,112,113,114,115,116,117,118,119,120,
				121,122,123,124,125,126,127,128,129,130,131,132,
				133,134,135,136,137,138,139,140,141,142,143,144,
				145,146,147,148,149,150,151,152,153,154,155,156,
				157,158,159,160,161,162,163,164,165,166,167,168,
				169,170,171,172,173,174,175,176,177,178,179,180,
				181,182,183,184,185,186,187,188,189,190,191,192,
				193,194,195,196,197,198,199,200,201,202,203,204,
				205,206,207,208,209,210,211,212,213,214,215,216,
				217,218,219,220,221,222,223,224,225,226,227,228,
				229,230,231,232,233,234,235,236,237,238,239,240;
	td=		1,2,3,4,5,6,7,8,9,10;
	tx=		1,2,3,4,5,6,7,8,9,10,
			11,12,13,14,15,16,17,18,19,20,
			21,22,23,24,25,26,27,28,29,30,
			31,32,33,34,35,36,37,38,39,40;
	ty=		1,2,3,4,5,6,7,8,9,10,
			11,12,13,14,15,16,17,18,19,20;
	tz=		1,2,3,4,5,6,7,8,9,10,
			11,12,13,14,15,16,17,18,19,20,
			21,22,23,24,25,26,27,28,29,30;
	txyz=		 	  1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12,
				 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24,
				 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36,
				 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48,
				 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60,
				 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72,
				 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84,
				 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96,
				 97, 98, 99,100,101,102,103,104,105,106,107,108,
				109,110,111,112,113,114,115,116,117,118,119,120,
				121,122,123,124,125,126,127,128,129,130,131,132,
				133,134,135,136,137,138,139,140,141,142,143,144,
				145,146,147,148,149,150,151,152,153,154,155,156,
				157,158,159,160,161,162,163,164,165,166,167,168,
				169,170,171,172,173,174,175,176,177,178,179,180,
				181,182,183,184,185,186,187,188,189,190,191,192,
				193,194,195,196,197,198,199,200,201,202,203,204,
				205,206,207,208,209,210,211,212,213,214,215,216,
				217,218,219,220,221,222,223,224,225,226,227,228,
				229,230,231,232,233,234,235,236,237,238,239,240;

//	three_double_dmn= 	 1, 2, 3, 4, 5, 6, 7, 8,
//				 9,10,11,12,13,14,15,16,
//				17,18,19,20,21,22,23,24,
//				-99,-99,-99,-99,-99,-99,-99,-99,
//				33,34,35,36,37,38,39,40,
//				41,42,43,44,45,46,47,48,
//				49,50,51,52,53,54,55,56,
//				-99,58,59,60,61,62,63,64,
//				65,66,67,68,69,70,71,72,
//				-99,74,75,76,77,78,79,-99,
//				1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5,
//				 9.5,10.5,11.5,12.5,13.5,14.5,15.5,16.5,
//				17.5,18.5,19.5,20.5,21.5,22.5,23.5,24.5,
//				-99.5,-99.5,-99.5,-99.5,-99.5,-99.5,-99.5,-99.5,
//				33.5,34.5,35.5,36.5,37.5,38.5,39.5,40.5,
//				41.5,42.5,43.5,44.5,45.5,46.5,47.5,48.5,
//				49.5,50.5,51.5,52.5,53.5,54.5,55.5,56.5,
//				-99.5,58.5,59.5,60.5,61.5,62.5,63.5,64.5,
//				65.5,66.5,67.5,68.5,69.5,70.5,71.5,72.5,
//				-99.5,74.5,75.5,76.5,77.5,78.5,79.5,-99.5;
				
	time_udunits = 876012, 876018, 876024;
	wnd_spd=		-999,0.5,1.5,0.5,1.5,0.5,1.5,0.5,
				0.5,-999,0.5,0.5,0.5,0.5,0.5,0.5,
				0.5,1.5,-999,1.5,0.5,1.5,0.5,1.5,
				0.5,0.5,0.5,-999,0.5,0.5,0.5,0.5,
  				1.5,1.5,1.5,1.5,-999,1.5,1.5,1.5,
				0.5,0.5,0.5,0.5,0.5,-999,0.5,0.5,
				2.5,2.5,2.5,2.5,2.5,2.5,-999,2.5,
				0.5,0.5,0.5,0.5,0.5,0.5,0.5,-999,
				0.5,0.5,0.5,0.5,0.5,0.5,0.5,0.5,
				0.5,0.5,2.5,0.5,0.5,2.5,0.5,0.5;
}







