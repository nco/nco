// -*-C++-*-
// Purpose: CDL file to generate netCDF4 test file for groups
// Created: 20110801 based on in.cdl

// Usage:
// NB: ncgen arguments depend on version:
// "-k netCDF-4" for netCDF >= 3.6.3, "-k hdf5" for netCDF < 3.6.3
// "-k netCDF-4 classic model" for netCDF >= 3.6.3, "-k hdf5-nc3" for netCDF < 3.6.3
// ncgen -k netCDF-4 -b -o ~/nco/data/in_grp.nc ~/nco/data/in_grp.cdl
// scp ~/nco/data/in_grp.cdl givre.ess.uci.edu:nco/data
// scp ~/nco/data/in_grp.nc dust.ess.uci.edu:/var/www/html/nco
// scp dust.ess.uci.edu:/var/www/html/nco/in_grp.nc ~/nco/data

// CDL Data constants:
// byte: 'a'
// char: "a"
// short: 1s
// int: 1 (no decimal point)
// float: 1.f (decimal point is required, f is required to distinguish from double)
// double: 1.0, 1.d, 1.0e-20 (decimal point is required, d is not required)
// CDL complex types:
// man ncgen describes all
// roulee:/data/zender/tmp/netcdf-4.2.1/nc_test/ref_tst_diskless2.cdl

// NCL usage:
// id_in=addfile("/home/zender/nco/data/in_grp.nc","r")
// print(id_in)
// list_filevars(id_in)
// ncks --get_file_info  ~/nco/data/in_grp.nc

netcdf in_grp {

 dimensions:
  lat=2;
  lev=3;
  lon=4;
  gds_crd=8;
  time=unlimited;
  tm2=unlimited;
  tm3=unlimited;
  vrt_nbr=2;
  
 variables:
  :Conventions = "CF-1.0";
  :history = "History global attribute.\n";
  :julian_day = 200000.04;
  :RCS_Header = "$Header: /data/zender/nco_20150216/nco/data/in_grp.cdl,v 1.62 2013-02-15 01:55:57 pvicente Exp $";
  float ilev(lev,vrt_nbr);
 ilev:purpose = "Cell boundaries for lev coordinate";
  double lat_gds(gds_crd);
 lat_gds:long_name = "Latitude";  
 lat_gds:standard_name = "latitude";
 lat_gds:units="degree";
 lat_gds:purpose = "1-D latitude coordinate referred to by geodesic grid variables";
  float lat(lat);
 lat:units = "degrees_north";
  float lev(lev);
 lev:units = "hybrid_sigma_pressure";
 lev:bounds = "ilev";
  float lon(lon);
 lon:units = "degrees_east";
  double lon_gds(gds_crd);
 lon_gds:long_name = "Longitude";
 lon_gds:standard_name = "longitude";
 lon_gds:units="degree";
 lon_gds:purpose = "1-D longitude coordinate referred to by geodesic grid variables";
  double time(time);
  float tm2(tm2);
 tm2:purpose = "a short record coordinate for testing mutiple record dimensions";
  float tm3(tm3);
 tm3:purpose = "another short record coordinate for testing mutiple record dimensions";
  float gds_crd(gds_crd);
 gds_crd:long_name = "Geodesic coordinate";
 gds_crd:units = "degree";
 gds_crd:purpose = "enumerated coordinate like those that might define points in a geodesic grid";
 gds_crd:coordinates = "lat_gds lon_gds";
  float scl;
  integer unique;
 unique:purpose = "the only variable of this name in this file, to test smallest possible access requests";    
  float area(lat);
 area:units = "meter2";
  float lat_lon(lat,lon);
  //float tm2_tm3(tm2,tm3);
  //tm2_tm3:purpose = "a variable containing mutiple record dimensions";
  //tm2_tm3:note = "ncdump prior to snapshot 20121116 and/or release netCDF 4.3 fails to print braces required to dis-ambiguate data sizes of mutiple record dimensions";
  //tm2_tm3:note2 = "ncgen from netCDF after ~201207 fails when ambiguous syntax (without braces) is used. Catch 22. Therefore remove tm2_tm3 from test file for now.";
  
 data:
  area=10.,10.;
  gds_crd=0,1,2,3,4,5,6,7;
  lat_gds=-90, -30,  -30,    0,   0, 30,  30,  90;
  lon_gds=  0,   0,  180,    0, 180,  0, 180,   0;
  lat=-90,90;
  lat_lon=1.,2.,3.,4.,5.,6.,7.,8;
  ilev=0,300,300,750,750,1013.25;
  lev=100,500,1000;
  lon=0,90,180,270;
  scl=1.0;
  time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
  tm2=1.,2.;
  tm3=1.,2.,3.;
  // 20130127: Braces are required to disambiguate correct record dimension sizes, but brace syntax but was not supported by ncgen until netCDF snapshots ~201211, i.e., post netCDF 4.2.1.1. Uggh.
  //tm2_tm3={1.,2.,3.},{4.,5.,6.};
  unique=73;
  //
  //g1
  //
 group: g1 { 
  variables:
    float lon(lon);
  lon:units = "g1 degrees_east";
    float scl;
    int g1v1;
    int v1;
  data:
    lon=0,90,180,270;
    scl=1.1;
    g1v1=1;
    v1=1;  
  group: g1g1 { 
    variables:
      float scl;
      int v1;
    data:
      scl=1.11;
      v1=11;
    } // end g1g1
  } // end g1
  
  //
  //g2
  //
 group: g2 { 
  variables:
    double time(time);
    float scl;
  data:
    time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
    scl=1.2;
  } // end g2
  
  //
  //g3
  //
 group: g3 {
  dimensions:
    rlev=3;
    time2=unlimited;
  variables:
    :g3_group_attribute = "g3_group_attribute";
    float rlev(rlev);
    rlev:purpose = "Monotonically decreasing coordinate pressure";
    double time2(time2);
    float rz(rlev);  
    float scl;
  data:
    time2=1.,2.;
    rz=0,5000,17000;
    scl=1.3;
    rlev=1000.,500.,100.;
    
  group: g3g1 {
    variables:
      float prs(rlev);
    prs:long_name="reverse pressure";
    data:
      prs=1.0,10.0,100.0;
    } // end g3g1
  } // end g3
  
  //
  //g4
  //
 group: g4 { 
  variables:
    int one_dmn_rec_var(time);
  one_dmn_rec_var:units = "second";
  data:
    one_dmn_rec_var=1,2,3,4,5,6,7,8,9,10;  
  } // end g4
  
  //
  //g5
  //
 group: g5 { // Level 1
  dimensions:
    rlev=3;
  variables:
    float rlev(rlev);
  data:
    rlev=10.,5.,1.;
  group: g5g1 { // Level 2
    variables:
      float rz(rlev);
    data:
      rz=1,2,3;
    } //end g6g1 
  } // end g5
  
  //
  //g6
  //
 group: g6 { // Level 1
  variables:
    float area(lat);
    float area1(lat);
  data:
    area=20.,30.;
    area1=21.,31.;
  group: g6g1 { // Level 2
    variables:
      float area(lat);
    data:
      area=40.,50.;
    } //end g6g1
  } // end g6
  
  //
  //g7
  //
 group: g7 { 
  dimensions:
    gds_crd=8;
  variables:
    float gds_crd(gds_crd);
  gds_crd:units = "degree";
  gds_crd:coordinates = "lat_gds lon_gds";
    float gds_var(gds_crd);
  gds_var:units = "meter";
  gds_var:coordinates = "lat_gds lon_gds";
    double lat_gds(gds_crd);
  lat_gds:units="degree";
    double lon_gds(gds_crd);
  lon_gds:units="degree";
  data:
    gds_crd=0,1,2,3,4,5,6,7;
    lat_gds=-90, -30,  -30,    0,   0, 30,  30,  90;
    lon_gds=  0,   0,  180,    0, 180,  0, 180,   0;
    gds_var=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8;
  } // end g7
  //
  //g8
  //
 group: g8 { 
  dimensions:
    lon=2,lev=3,vrt_nbr=2;
  variables:
    float lev(lev);
    float lon(lon);
    lev:units = "hybrid_sigma_pressure";
    lev:bounds = "ilev";
    float vrt_nbr(vrt_nbr);
    float ilev(lev,vrt_nbr);
  data:
    lon=-180,0; 
    lev=100,500,1000;
    ilev=0,300,300,750,750,1013.25;
    vrt_nbr=1,2;
  } // end g8
  
  //
  //g9
  //
 group: g9 { // Level 1
  group: g9g1 { // Level 2
    variables:
      int v6;
    data:
      v6=63;
    group: g9g1g1 { // Level 3
      group: g9g1g1g1 { // Level 4
	  :mtd_grp = "Group metadata from g9g1g1g1, a group with no variables, to test whether group metadata are copied to ancestor groups of extracted variables";
	group: g9g1g1g1g1 { // Level 5
	  group: g9g1g1g1g1g1 { // Level 6
	    group: g9g1g1g1g1g1g1 { // Level 7
	      variables:
		int v7;
	      data:
		v7=73;
	      } // end g9g1g1g1g1g1g1
	    } // end g9g1g1g1g1g1
	  } // end g9g1g1g1g1
	} // end g9g1g1g1
      } // end g9g1g1
    } // end g9g1
  } // end g9

 group: g10 { // Level 1
  variables:
    float two_dmn_rec_var(time,lev);
    float three_dmn_rec_var(time,lat,lon);
  data:
    two_dmn_rec_var=1.,2.0,3.,
      1.,2.1,3.,
      1.,2.2,3.,
      1.,2.3,3.,
      1.,2.4,3.,
      1.,2.5,3.,
      1.,2.6,3.,
      1.,2.7,3.,
      1.,2.8,3.,
      1.,2.9,3.;
    three_dmn_rec_var= 	 1, 2, 3, 4, 5, 6, 7, 8,
      9,10,11,12,13,14,15,16,
      17,18,19,20,21,22,23,24,
      25,26,27,28,29,30,31,32,
      33,34,35,36,37,38,39,40,
      41,42,43,44,45,46,47,48,
      49,50,51,52,53,54,55,56,
      57,58,59,60,61,62,63,64,
      65,66,67,68,69,70,71,72,
      73,74,75,76,77,78,79,80;
  } // end g10

 group: g11 { // Level 1
    // Purpose: Test netCDF4-specific atomic types
  variables:
    int64 int64_var;
  int64_var:long_name = "int64-type variable";
    
    string string_var;
  string_var:long_name = "string-type variable";
    
    ubyte ubyte_var;
  ubyte_var:long_name = "ubyte-type variable";
    
    uint uint_var;
  uint_var:long_name = "uint-type variable";
    
    uint uint_arr(lat);
  uint_arr:long_name = "uint-type array variable";
    
    uint64 uint64_var;
  uint64_var:long_name = "uint64-type variable";
    
    ushort ushort_var;
  ushort_var:long_name = "ushort-type variable";
  data:
    int64_var=9223372036854775807; // LLONG_MAX = 9223372036854775807, NC_FILL_INT64 is -9223372036854775806LL
    string_var="If you prick us, do we not bleed? If you tickle us, do we not laugh? If you poison us, do we not die? And if you wrong us, shall we not revenge?";
    ubyte_var='z'; // UCHAR_MAX = 255, NC_FILL_UBYTE = 255
    // 20130208: netCDF 4.2.1 and snapshots to date fail as nc_get_var1_uint() returns -60 = NetCDF: Numeric conversion not representable on following (valid) input value. Works for 0, though, and for arrays.
    // uint_var=4294967295; // UINT_MAX = 4294967295, NC_FILL_UINT is 4294967295U
    uint_var=0; // UINT_MAX = 4294967295, NC_FILL_UINT is 4294967295U
    uint_arr=4294967295,4294967295; // UINT_MAX = 4294967295, NC_FILL_UINT is 4294967295U
    uint64_var=18446744073709551615; // ULLONG_MAX = 18446744073709551615, NC_FILL_UINT is 18446744073709551614ULL
    ushort_var=65535; // USHRT_MAX = 65535, NC_FILL_USHORT = 65535
 } // end g11

 group: g12 { // Level 1
    // Purpose: Test netCDF4 vlen type
    // 20130208: ncgen from netCDF 4.2.1- broken for vlen types
    // Probably broken on all snapshots until ~201211 because brace-handling broken
  types:
    int(*) vlen_t;
  variables:
    vlen_t vlen_var;
  data:
    vlen_var={17,18,19};
  } // end g12

 group: g13 { // Level 1
    // Purpose: Test netCDF4 opaque type
  types:
    opaque(11) opaque_t;
  } // end g13

 group: g14 { // Level 1
    // Purpose: Test netCDF4 enum type
  types:
    ubyte enum enum_t {Clear=0,Cumulonimbus=1,Stratus=2};
  variables:
    enum_t cloud_flg(lon);
  data:
    cloud_flg=Stratus,Stratus,Cumulonimbus;
  } // end g14

 group: g15 { // Level 1
    // Purpose: Test netCDF4 compound type
  types:
    compound cmpd_t {vlen_t f1;enum_t f2;};
  variables:
    cmpd_t compound_var;
  data:
    compound_var={{3,4,5},Stratus};
  } // end g15
  
  
  //
  //g16 
  //
  // Test variables and dimensions in and out of scope
  // Use case of variable in scope of dimension:
  // dimension /lon 
  // variable /g1/lon(lon)
  // Use case of variable NOT in scope of dimension:
  // variable /lon
  // dimension /g1/lon
  //
  // Test dimensions with no associated coordinate variable
  //
  group: g16 { 
    dimensions:
    lon1=4;  //dimension that has a coordinate variable down in scope at /g16/g16g1/lon1(lon1)
    lon2=4;  //dimension that does NOT have a coordinate variable anywhere 
    variables:
    float lat1(lat);
    //NOTE: attempting to define float lat1(lat1); is not legal: ncgen: Undefined or forward referenced dimension: lat1
    //But we can try to define a dimension lat1 anyway down in the group path for NCO testing/sanity check
    float lon2_var(lon2); //variable with no associated coordinate variable
    data:
    lat1=1.,2.;
    lon2_var=1.,2.,3.,4.; 
    
    group: g16g1 { 
     dimensions:
     lat1=2; //dimension that has a variable /lat1 down in *illegal* scope 
     variables:
     float lon1(lon1);  //coordinate variable /g16/g16g1/lon1(lon1) that has dimension /lon1 in scope
     float lon1_var(lon1); //variable with  associated coordinate variable down in scope at /lon1
     data:
     lon1=1.,2.,3.,4.;
     lon1_var=1.,2.,3.,4.; 
      } // end g16g1 
  } // end g16
  
  

} // end root group
