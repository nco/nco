// Generate netCDF file with:
// ncgen -k netCDF-4 -b -o ~/nco/data/cmip5.nc ~/nco/data/cmip5.cdl

netcdf cmip5 {
  dimensions:
  time=unlimited;
 
  //
  //cesm
  //
  group: cesm { 
  variables:
  float tas(time);
  data:
  tas=0,0,0,0;
  } // end cesm
  
  //
  //ecmwf
  //
  group: ecmwf { 
  variables:
  float tas(time);
  data:
  tas=1,1,1,1;
  } // end ecmwf
  
  //
  //gfdl
  //
  group: gfdl { 
  variables:
  float tas(time);
  data:
  tas=2,2,2,2;
  } // end gfdl

} // end root group
