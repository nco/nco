// Purpose: CDL file to generate netCDF test file

// Usage:
// ncgen -b -o in.nc in.cdl
// ncgen -b -o ${HOME}/nco/data/in.nc ${HOME}/nco/data/in.cdl
// mswrite -t 365 ~/nco/data/in.nc /ZENDER/tmp/in.nc
// mswrite -t 365 ~/nco/data/in.nc /ZENDER/tmp/h0001.nc
// mswrite -t 365 ~/nco/data/in.nc /ZENDER/tmp/h0002.nc
// mswrite -t 365 ~/nco/data/in.nc /ZENDER/tmp/h0003.nc
// mswrite -t 365 ~/nco/data/in.nc /ZENDER/tmp/h0004.nc
// msrcp -period 365 ~/nco/data/in.nc mss:/ZENDER/tmp/in.nc
// msrcp -period 365 ~/nco/data/in.nc mss:/ZENDER/tmp/h0001.nc
// msrcp -period 365 ~/nco/data/in.nc mss:/ZENDER/tmp/h0002.nc
// msrcp -period 365 ~/nco/data/in.nc mss:/ZENDER/tmp/h0003.nc
// msrcp -period 365 ~/nco/data/in.nc mss:/ZENDER/tmp/h0004.nc

// WARNING: Changing values of variables below, especially coordinate variables, will affect the outcome of nco_tst.sh test script
// Other programs, e.g., ~/f/fff.F90, ~/c++/ccc.cc, ~/c/c.c may also break
// In particular, do not change the number of elements in the record coordinate, time, without simultaneously changing the number of data in all the record variables

// Data constants in CDL:
// byte: 'a'
// char: "a"
// short: 1s
// int: 1 (no decimal point)
// float: 1.f (decimal point is required, f is required to distinguish from double)
// double: 1.0, 1.d, 1.0e-20 (decimal point is required, d is not required)

// NCL usage:
// id_in=addfile("/home/zender/nco/data/in.nc","r")
// print(id_in)
// list_filevars(id_in)

netcdf in {
dimensions:
	bnd=2,lat=2,lev=3,rlev=3,lon=4,char_dmn_lng=80,char_dmn_sml=4,fl_dim=3,lsmlev=6,wvl=2,time=unlimited;
variables:
	:Conventions = "NCAR-CSM";
	:history = "History global attribute.\n";
	:julian_day = 200000.04;
	:RCS_Header = "$Header: /data/zender/nco_20150216/nco/data/in.cdl,v 1.38 2002-08-21 11:47:41 zender Exp $";

	float lat(lat);
	float lat_var(lat);
	float lat_wgt(lat);
	float lev(lev);
	lev:purpose = "Monotonically increasing coordinate pressure";
	lev:units = "hybrid_sigma_pressure";
	lev:positive = "down";
	lev:A_var = "hyam";
	lev:B_var = "hybm";
	lev:P0_var = "P0";
	lev:PS_var = "PS";
	lev:bounds = "ilev";
	float rlev(rlev);
	rlev:purpose = "Monotonically decreasing coordinate pressure";
	float lon(lon);
	double time(time);
	float lsmlev(lsmlev);
	lsmlev:purpose = "Homebrew level coordinate for LSM";
	lsmlev:long_name = "Soil depth";
	lsmlev:units = "meter";
	float wvl(wvl);
	wvl:long_name = "Wavelength";
	wvl:units = "meter";

	float hyam(lev);
	hyam:long_name = "hybrid A coefficient at layer midpoints";

	float hybm(lev);
	hybm:long_name = "hybrid B coefficient at layer midpoints";

	float P0;
	P0:long_name = "reference pressure";
	P0:units = "pascal";

	float PS(time,lat,lon);
	PS:long_name = "surface pressure";
	PS:units = "pascal";

	char fl_dim(fl_dim);
	fl_dim:long_name = "Character coordinate";
	fl_dim:units = "[chr]";

	int nbdate;
	nbdate:long_name = "base date as 6 or 8 digit integer (YYMMDD or YYYYMMDD)";
	int date(time);
	date:long_name = "current date as 6 or 8 digit integer (YYMMDD or YYYYMMDD)";

	float lon_wgt(lon);
	lon_wgt:long_name = "Gaussian weights";
	lon_wgt:purpose = "Gaussian weights which sum to two for n = 4. These weights are all have floor of 0.0 so should cause SIGFPE when applied to integer types in weighted average.";

	float msk_prt_mss_prt(lon);
	msk_prt_mss_prt:long_name = "partial mask, partial missing value example";
	msk_prt_mss_prt:missing_value = 1.0e36f;

	float mss_val(lon);
	mss_val:long_name = "partial missing value example";
	mss_val:missing_value = 1.0e36f;

	float fll_val(lon);
	fll_val:long_name = "_FillValue example";
	fll_val:_FillValue = -999.0f;

	float no_mss_val(lon);
	no_mss_val:long_name = "no missing value";

	float val_one_mss(lat);
	val_one_mss:long_name = "one regular value, one missing value";
	val_one_mss:missing_value = 1.0e36f;

	short pck;
	pck:long_name = "Packed scalar variable";
	pck:note = "Packed value is 1s, unpacked is 2.0d0*1s + 1.0d0 = 3.0d0.";
	pck:scale_factor = 2.0d;
	pck:add_offset = 1.0d;

	short pck_arr(lon);
	pck_arr:long_name = "Packed array";
	pck_arr:note = "Packed value is -32767s, 0s, 1s, 32767s, unpacked is same in double";
	pck_arr:scale_factor = 1.0d;
	pck_arr:add_offset = 0.0d;

	double upk;
	upk:long_name = "Unpacked scalar variable";
	upk:note = "Unpacked value is 3.0d0, upk=unpack(pck)= 2.0d0*1s + 1.0d0 = 3.0d0. Packing this variable should create an NC_SHORT scalar = 0s with packing attribute add_offset=3.0d";

	double upk_arr(lon);
	upk_arr:long_name = "Unpacked array";
	upk_arr:note = "Unpacked value is -32767.d, 0.d, 1.d, 32767.d, packed is same in short. Packing algorithm should yield an NC_SHORT array = [] with packing attributes scale_factor=1.0d, add_offset=0.0d";

	int val_one_int;
	val_one_int:long_name = "scalar equal to 1";
	val_one_int:missing_value = -99l;

	int val_one_one_int(lat);
	val_one_one_int:long_name = "1, 1";
	val_one_one_int:missing_value = -99l;

	short val_max_max_sht(lat);
	val_max_max_sht:long_name = "17000, 17000";
	val_max_max_sht:missing_value = -99s;

	int val_one_mss_int(lat);
	val_one_mss_int:long_name = "1, mss_val";
	val_one_mss_int:missing_value = -99l;

	float val_half;
	val_half:long_name = "Scalar with value 0.5";
	val_half:missing_value = 1.0e36f;

	float val_half_half(lat);
	val_half_half:long_name = "0.5,0.5";
	val_half_half:missing_value = 1.0e36f;

	float wgt_one(lat);
	wgt_one:long_name = "all values are one";

	float mss_val_all(lon);
	mss_val_all:long_name = "all missing values example";
	mss_val_all:missing_value = 1.0e36f;

	float scalar_var;
	scalar_var:long_name = "scalar variable";
	scalar_var:units = "Fraction";

	float float_var;
	float_var:long_name = "float";

	double double_var;
	double_var:long_name = "double";

	int int_var;
	int_var:long_name = "int";

	short short_var;
	short_var:long_name = "short";

	char char_var;
	char_var:long_name = "char";

	char char_var_space;
	char_var_space:long_name = "Character variable with whitespace on ends";

	char char_var_nul;
	char_var_nul:long_name = "Character variable containing one NUL";

	char char_var_multinul(lev);
	char_var_multinul:long_name = "Character variable containing multiple NULs";

	char fl_nm(char_dmn_lng);
	fl_nm:long_name = "Variable contains a file name";

	char fl_nm_arr(fl_dim,char_dmn_lng);
	fl_nm_arr:long_name = "Variable that contains a short array of file names";
	fl_nm_arr:units = "[sng]";

	char non_nul_trm_char_one_dim(char_dmn_sml);
	non_nul_trm_char_one_dim:long_name = "Variable contains a one-dimensional array of characters that is not NUL-terminated";
	non_nul_trm_char_one_dim:units = "[chr]";

	char non_nul_trm_char_two_dim(fl_dim,char_dmn_sml);
	non_nul_trm_char_two_dim:long_name = "Variable contains a two-dimensional array of characters that are not NUL-terminated";
	non_nul_trm_char_two_dim:units = "[chr]";

	byte byte_var;
	byte_var:long_name = "byte";

	float zero;
	zero:long_name = "zero";

	float one;
	one:long_name = "one";

	float two;
	two:long_name = "two";

	float three;
	three:long_name = "three";

	float four;
	four:long_name = "four";

	float negative_one;
	negative_one:long_name = "negative one";

	float lev_var(lev);
	lev_var:long_name = "lev_var";

	float lev_wgt(lev);
	lev_wgt:long_name = "lev_wgt";

	float g;
	g:long_name = "g";

	float z(lev);
	z:long_name = "Height";
	z:units = "meter";
	z:purpose = "Height stored with a monotonically increasing coordinate";

	float rz(rlev);
	rz:long_name = "Height";
	rz:units = "meter";
	rz:purpose = "Height stored with a monotonically decreasing coordinate";

	float one_dmn_var(bnd);

	float att_var;
	att_var:byte_att = '\0';
	att_var:char_att = "Sentence one.\nSentence two.\n";
	att_var:short_att = 37s;
	att_var:int_att = 73l;
	att_var:float_att = 73.0f,72.0f,71.0f;
	att_var:double_att = 73.0d;

	int bnd_var(lev,bnd);
	bnd_var:byte_att = '\0';
	bnd_var:char_att = "Sentence one.\nSentence two.\n";
	bnd_var:short_att = 37s;
	bnd_var:int_att = 73;
	bnd_var:float_att = 73.f;
	bnd_var:double_att = 73.d;

	float three_dmn_var(lat,lev,lon);
	three_dmn_var:long_name = "three dimensional variable with CCM coordinate convention C=[lat,lev,lon], Fortran=(lon,lev,lat)";
	three_dmn_var:units = "Fraction";

	float three_dmn_var_crd(lev,lat,lon);
	three_dmn_var_crd:long_name = "three dimensional variable with COORDS coordinate convention C=[lev,lat,lon], Fortran=(lon,lat,lev)";
	three_dmn_var_crd:units = "Fraction";

	float prs_sfc(time,lat,lon);
	prs_sfc:long_name = "Surface pressure";
	prs_sfc:units = "pascal";

	float two_dmn_var(lat,lev);
	two_dmn_var:long_name = "two dimensional variable";
	two_dmn_var:units = "Fraction";

	float mask(lat,lon);
	mask:long_name = "mask variable like ORO";
	mask:units = "Fraction";

	float ORO(lat,lon);
	ORO:long_name = "Orography";
	ORO:units = "Fraction";

	float weight(lat);
	weight:long_name = "Gaussian weight";
	weight:units = "Fraction";

	float gw(lat);
	gw:long_name = "gw variable like gw";
	gw:units = "Fraction";

	float rec_var_flt(time);
	rec_var_flt:long_name = "record variable, float";

	double rec_var_dbl(time);
	rec_var_dbl:long_name = "record variable, double";

	int one_dmn_rec_var(time);
	one_dmn_rec_var:long_name = "one dimensional record variable";
	one_dmn_rec_var:units = "second";

	float tpt(time);
	tpt:long_name = "Temperature";
	tpt:units = "kelvin";

	double rec_var_dbl_mss_val_dbl_upk(time);
	rec_var_dbl_mss_val_dbl_upk:long_name = "record variable, double, with double missing values";
	rec_var_dbl_mss_val_dbl_upk:purpose = "This variable is used to generate the packed variable rec_var_dbl_mss_val_dbl_pck, so its missing_value should not be too far out of range, i.e., it should be representable by a short";
	rec_var_dbl_mss_val_dbl_upk:missing_value = -999.;

	short rec_var_dbl_mss_val_dbl_pck(time);
	rec_var_dbl_mss_val_dbl_pck:long_name = "record variable, double, with double missing values, packed";
	rec_var_dbl_mss_val_dbl_pck:purpose = "Packed version of rec_var_dbl_mss_val_dbl_upk";
	rec_var_dbl_mss_val_dbl_pck:missing_value = -999s;
        rec_var_dbl_mss_val_dbl_pck:scale_factor = -9.15541313801785e-05 ;
        rec_var_dbl_mss_val_dbl_pck:add_offset = 5. ;

	float rec_var_flt_mss_val_flt(time);
	rec_var_flt_mss_val_flt:long_name = "record variable, float, with float missing values";
	rec_var_flt_mss_val_flt:missing_value = 1.0e36f;

	float rec_var_flt_mss_val_dbl(time);
	rec_var_flt_mss_val_dbl:long_name = "record variable, float, with double missing values";
	rec_var_flt_mss_val_dbl:missing_value = 1.0e36d;

	float rec_var_flt_mss_val_int(time);
	rec_var_flt_mss_val_int:long_name = "record variable, float, with integer missing values";
	rec_var_flt_mss_val_int:missing_value = -999;

	int rec_var_int_mss_val_int(time);
	rec_var_int_mss_val_int:long_name = "record variable, integer, with integer missing values";
	rec_var_int_mss_val_int:missing_value = -999;

	int rec_var_int_mss_val_flt(time);
	rec_var_int_mss_val_flt:long_name = "record variable, integer, with float missing values";
	rec_var_int_mss_val_flt:missing_value = -999.0f;

	int rec_var_int_mss_val_dbl(time);
	rec_var_int_mss_val_dbl:long_name = "record variable, integer, with double missing values";
	rec_var_int_mss_val_dbl:missing_value = -999.0;

	int rec_var_dbl_mss_val_dbl_pck_lng(time);
	rec_var_dbl_mss_val_dbl_pck_lng:long_name = "record variable, double packed as long, with double missing values";
	rec_var_dbl_mss_val_dbl_pck_lng:purpose = "although not usual, packing doubles into longs (rather than shorts) is still a considerable cost savings";
	rec_var_dbl_mss_val_dbl_pck_lng:missing_value = -999;
        rec_var_dbl_mss_val_dbl_pck_lng:scale_factor = -9.15541313801785e-05 ;
        rec_var_dbl_mss_val_dbl_pck_lng:add_offset = 5. ;

	char one_dmn_rec_var_sng(time);
	one_dmn_rec_var_sng:long_name = "one dimensional record variable of string";

	float time_lon(time,lon);
	time_lon:long_name = "Record variable of longitude coordinate";

	char two_dmn_rec_var_sng(time,lev);
	two_dmn_rec_var_sng:long_name = "two dimensional record variable of string";

	float two_dmn_rec_var(time,lev);
	two_dmn_rec_var:long_name = "two dimensional record variable";
	two_dmn_rec_var:units = "watt meter-2";

	float three_dmn_rec_var(time,lat,lon);
	three_dmn_rec_var:long_name = "three dimensional record variable";
	three_dmn_rec_var:units = "watt meter-2";

	double three_dmn_var_dbl(time,lat,lon);
	three_dmn_var_dbl:long_name = "three dimensional record variable of type double";
	three_dmn_var_dbl:units = "watt meter-2";
	three_dmn_var_dbl:missing_value = -99 ;

	int three_dmn_var_int(time,lat,lon);
	three_dmn_var_int:long_name = "three dimensional record variable of type int";
	three_dmn_var_int:units = "watt meter-2";
	three_dmn_var_int:missing_value = -99 ;
	
	short three_dmn_var_sht(time,lat,lon);
	three_dmn_var_sht:long_name = "three dimensional record variable";
	three_dmn_var_sht:units = "watt meter-2";
	three_dmn_var_sht:missing_value = -99 ;

	float four_dmn_rec_var(time,lat,lev,lon);
	four_dmn_rec_var:long_name = "four dimensional record variable";
	four_dmn_rec_var:units = "watt meter-2";

data:
	ORO=1.,1.,1.,1.,1.,1.,1.,1.;
	att_var=10.;
	bnd_var=1,2,3,4,5,6;
	byte_var='z';
	char_var="z";
	char_var_multinul="\b\n\0";
	char_var_nul='\0';
	char_var_space=" ";
	double_var=10.;
	fl_dim="a","b","3";
	fl_nm="/home/zender/nco/data/in.cdl";
	float_var=10.;
	g=9.8;
	gw=10.,10.;
	hyam=0.0802583,0.0438226,0.0;
	hybm=0.0187849,0.457453,0.992528;
	P0=100000;
	lat=-90,90;
	lat_var=1.,2.;
	lat_wgt=1.,2.;
	lsmlev=0.05,0.1,0.2,0.5,1.0,3.0;
	lev=100,500,1000;
	lev_var=100.,500.,1000.;
	lev_wgt=10,2,1;
	lon=0,90,180,270;
	lon_wgt=0.347855,0.652145,0.652145,0.347855;
	mask=0.,1.,0.,0.,1.,1.,0.,2.;
//	mask=0.,0.,0.,0.,0.,0.,0.,0.;
//	mask=1.,1.,1.,1.,1.,1.,1.,1.;
	fll_val=73,-999,73,-999;
	msk_prt_mss_prt=0.5,1.0e36,1.5,1.0e36;
	mss_val=73,1.0e36,73,1.0e36;
	mss_val_all=1.0e36,1.0e36,1.0e36,1.0e36;
	negative_one=-1.;
	no_mss_val=73,1.0e36,73,1.0e36;
	non_nul_trm_char_one_dim='a','b';
	non_nul_trm_char_two_dim="abcd","efgh","ijkm";
	one=1.;
	four=4.;
	one_dmn_rec_var=1,2,3,4,5,6,7,8,9,10;
	one_dmn_rec_var_sng="Hello Wor";
	one_dmn_var=1.,10.;
	pck=1;
	pck_arr=-32767,0,1,32767;
	upk=3.;
	upk_arr=-32767.,0.,1.,32767.;
	rec_var_dbl=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	rec_var_flt=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	rec_var_dbl_mss_val_dbl_pck=-999,32767,21845,10922,0,-10922,-21845,-32767,-999,-999;
	rec_var_dbl_mss_val_dbl_upk=-999.,2.,3.,4.,5.,6.,7.,8.,-999.,-999.;
	rec_var_flt_mss_val_dbl=1.0e36,2.,3.,4.,5.,6.,7.,8.,1.0e36,1.0e36;
	rec_var_flt_mss_val_flt=1.0e36,2.,3.,4.,5.,6.,7.,8.,1.0e36,1.0e36;
	rec_var_flt_mss_val_int=-999.,2.,3.,4.,5.,6.,7.,8.,-999.,-999.;
	rec_var_int_mss_val_int=-999,2,3,4,5,6,7,8,-999,-999;
	rec_var_int_mss_val_flt=-999,2,3,4,5,6,7,8,-999,-999;
	rec_var_dbl_mss_val_dbl_pck_lng=-999,32767,21845,10922,0,-10922,-21845,-32767,-999,-999;
	rec_var_int_mss_val_dbl=-999,2,3,4,5,6,7,8,-999,-999;
	rlev=1000,500,100;
	rz=0,5000,17000;
	scalar_var=10.;
	short_var=10;
	three=3.;
	three_dmn_var=0.,1.,2.,3.,4.,5.,6.,7.,8.,9.,10.,11.,12.,13.,14.,15.,16.,17.,18.,19.,20.,21.,22.,23.;
	three_dmn_var_crd=0.,1.,2.,3.,12.,13.,14.,15.,4.,5.,6.,7.,16.,17.,18.,19.,8.,9.,10.,11.,20.,21.,22.,23.;
	time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	tpt=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8,273.9,273.10;
	two=2.;
	two_dmn_var=1.5,5.5,9.5,13.5,17.5,21.5;
	val_half=0.5;
	val_half_half=0.5,0.5;
	val_max_max_sht=17000,17000;
	val_one_int=1;
	val_one_mss=1.,1.0e36;
	val_one_mss_int=1,-99;
	val_one_one_int=1,1;
	weight=10.,10.;
	wgt_one=1.,1.;
	wvl=0.5e-6,1.0e-6;
	z=17000,5000,0;
	zero=0.;
 	date=640312,640313,640314,640315,640316,640317,640318,640319,640320,640321;
 	int_var=10;
 	nbdate=640312;
	fl_nm_arr="/data/zender/dstccm04/dstccm04_8589_01.nc",
		"/data/zender/dstccm04/dstccm04_8589_02.nc",
		"/data/zender/dstccm04/dstccm04_8589_03.nc";
	time_lon=0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0;
	two_dmn_rec_var_sng="abc",
				"bcd",
				"cde",
				"def",
				"efg",
				"fgh",
				"ghi",
				"hij",
				"jkl",
				"klm";
	two_dmn_rec_var=1.,2.0,3.,
			1.,2.1,3.,
			1.,2.2,3.,
			1.,2.3,3.,
			1.,2.4,3.,
			1.,2.5,3.,
			1.,2.6,3.,
			1.,2.7,3.,
			1.,2.8,3.,
			1.,2.9,3.;
	three_dmn_rec_var= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
  				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				73,74,75,76,77,78,79,80;
	prs_sfc=		 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
  				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				73,74,75,76,77,78,79,80;
	PS=			101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
  				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325;
	three_dmn_var_dbl= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				-99,-99,-99,-99,-99,-99,-99,-99,
				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				-99,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				-99,74,75,76,77,78,79,-99;
	three_dmn_var_int= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				-99,-99,-99,-99,-99,-99,-99,-99,
				25,26,27,28,29,30,31,32,
				33,34,35,36,37,38,39,40,
				41,-99,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				-99,58,59,60,-99,62,63,64,
				65,-99,67,68,69,70,71,72,
				-99,74,75,-99,77,78,79,80;
	three_dmn_var_sht= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 -99,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
				-99,34,35,-99,37,38,39,40,
				41,42,43,44,-99,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,-99,61,62,63,64,
				65,66,67,68,69,70,71,72,
				-99,-99,-99,-99,-99,-99,-99,-99;

	four_dmn_rec_var= 	  1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12,
				 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24,
				 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36,
				 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48,
				 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60,
				 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72,
				 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84,
				 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96,
				 97, 98, 99,100,101,102,103,104,105,106,107,108,
				109,110,111,112,113,114,115,116,117,118,119,120,
				121,122,123,124,125,126,127,128,129,130,131,132,
				133,134,135,136,137,138,139,140,141,142,143,144,
				145,146,147,148,149,150,151,152,153,154,155,156,
				157,158,159,160,161,162,163,164,165,166,167,168,
				169,170,171,172,173,174,175,176,177,178,179,180,
				181,182,183,184,185,186,187,188,189,190,191,192,
				193,194,195,196,197,198,199,200,201,202,203,204,
				205,206,207,208,209,210,211,212,213,214,215,216,
				217,218,219,220,221,222,223,224,225,226,227,228,
				229,230,231,232,233,234,235,236,237,238,239,240;
}







