// -*-C++-*-

// Purpose: CDL file to generate NCZarr-compatible test file with netCDF4 atomic types for NCO
// Derived by removing NCZarr incompatibilities from in.cdl
// Changes include:
// 1. Change time from NC_UNLIMITED to fixed size 10
// 2. Add netCDF4 types from in_4.cdl
// 3. Remove all variables and attributes of string type
// 4. Make all scalars use degenerate (size = 1) "scalar" dimension as (hopefully) temporary workaround to https://github.com/Unidata/netcdf-c/issues/2485
// 5. 20220827: Eliminate Lat,Lon dimensions 
// 6. 20220830: Restore variables/attributes of string type after PR #2492 by D. Heimbigner added support for strings
// 7. Report regressions in string handling to Unidata
// 8. 20220906 Re-test variables/attributes of string type after PR #2497 by D. Heimbigner fixed support for strings. Strings now work as advertised
// 9. 20220907 Report "Unmatched untrace: fcn=ncz_get_var_meta expected=NCZ_inq_var_filter_info" issue
// 10. Remove degenerate "scalar" dimension which NCZarr now supports
// 11. Restore NC_UNLIMITED after PR #2744 by D. Heimbigner added support for unlimited dimensions
// 12. Temporarily eliminate NC_UNLIMITED dimension so NCO 5.1.9+ distribution does not break when building with netCDF <= 4.9.2

// Usage:
// netCDF4: ncgen arguments depend on version:
// "-k netCDF-4" for netCDF >= 3.6.3, "-k hdf5" for netCDF < 3.6.3
// "-k netCDF-4 classic model" for netCDF >= 3.6.3, "-k hdf5-nc3" for netCDF < 3.6.3
// ncgen -k netCDF-4 -b -o in_zarr4.nc in_zarr4.cdl
// ncgen -k netCDF-4 -b -o ${HOME}/nco/data/in_zarr4.nc ${HOME}/nco/data/in_zarr4.cdl
// ncgen -lb -o "file://${HOME}/in_zarr4#mode=nczarr,file" ${HOME}/nco/data/in_zarr4.cdl
// ncks -O -4 "file://${HOME}/in_zarr4#mode=nczarr,file" ~/in_zarr4.nc

// URL:
// http://dust.ess.uci.edu/nco/in_zarr4.nc
// http://dust.ess.uci.edu/nco/in_zarr4.nc
// http://thredds-test.ucar.edu/thredds/dodsC/testdods/in_zarr4.nc

// netCDF3:
// ncgen -b -o in_zarr4.nc in_zarr4.cdl
// ncgen -b -o ${HOME}/nco/data/in_zarr4.nc ${HOME}/nco/data/in_zarr4.cdl
// scp ~/nco/data/in_zarr4.cdl ~/nco/data/in_4.nc dust.ess.uci.edu:nco/data
// scp ~/nco/data/in_zarr4.nc ~/nco/data/in_4.nc dust.ess.uci.edu:/var/www/html/nco
// scp ~/nco/data/in_zarr4.nc ~/nco/data/in_4.nc dust.ess.uci.edu:/var/www/html/dodsdata
// mswrite -t 365 ~/nco/data/in_zarr4.nc /ZENDER/tmp/in_zarr4.nc
// mswrite -t 365 ~/nco/data/in_zarr4.nc /ZENDER/tmp/h0001.nc
// mswrite -t 365 ~/nco/data/in_zarr4.nc /ZENDER/tmp/h0002.nc
// mswrite -t 365 ~/nco/data/in_zarr4.nc /ZENDER/tmp/h0003.nc
// mswrite -t 365 ~/nco/data/in_zarr4.nc /ZENDER/tmp/h0004.nc
// msrcp -period 365 ~/nco/data/in_zarr4.nc mss:/ZENDER/tmp/in_zarr4.nc
// msrcp -period 365 ~/nco/data/in_zarr4.nc mss:/ZENDER/tmp/h0001.nc
// msrcp -period 365 ~/nco/data/in_zarr4.nc mss:/ZENDER/tmp/h0002.nc
// msrcp -period 365 ~/nco/data/in_zarr4.nc mss:/ZENDER/tmp/h0003.nc
// msrcp -period 365 ~/nco/data/in_zarr4.nc mss:/ZENDER/tmp/h0004.nc

// WARNING: Changing values of variables below, especially coordinate variables, affects outcome of nco_tst.pl test script
// Other programs, e.g., ~/f/fff.F90, ~/c++/ccc.cc, ~/c/c.c may also break
// In particular, do not change number of elements in record coordinate, time, without simultaneously changing number of data in all record variables
// My (and NCO's) convention is that the _FillValue, if any, of any packed variable should be of the same type as the expanded variable. Hence _FillValue, add_offset, and scale_factor should all be of the same type. Variables that do not adhere to this convention are not supported.

// Bugs:
// Some triggering bugs were moved to buggy.cdl to prevent non-builds
// ncgen 4.0.0--4.3.2 crashes on 'l' or 'L' syntax when generating netCDF4-classic (but not netCDF3 or netCDF4) files until 20141010 (NCF-318)

// CDL Data constants:
// http://www.unidata.ucar.edu/software/netcdf/docs/netcdf/CDL-Syntax.html
// byte: 'a'
// char: "a"
// short: 1s
// int: 1 (no decimal point)
// long: 1 (_not_ 1l;) (long is synonym for int in netCDF3)
// float: 1.f (decimal point is required, f is required to distinguish from double)
// double: 1.0, 1.d, 1.0e-20 (decimal point is required, d is not required)
// CDL complex types:
// roulee:/data/zender/tmp/netcdf-4.2.1/nc_test/ref_tst_diskless2.cdl

// NCL usage:
// id_in=addfile("/home/zender/nco/data/in.nc","r")
// print(id_in)
// list_filevars(id_in)

netcdf in_zarr4 {
dimensions:
//dgn=1,bnd=2,lat=2,lat_grd=3,lev=3,rlev=3,ilev=4,lon=4,lon_grd=5,char_dmn_lng80=80,char_dmn_lng26=26,char_dmn_lng04=4,date_dmn=5,fl_dmn=3,lsmlev=6,wvl=2,time_int_udunits=1;time_udunits=3;lon_T42=128,lat_T42=64,lat_times_lon=8,gds_crd=8,gds_ncd=8,lon_cal=10,lat_cal=10,Lon=4,Lat=2,pck_crd=4,vrt_nbr=2,time=10;
// 20220827: Eliminate Lat,Lon dimensions
//dgn=1,bnd=2,lat=2,lat_grd=3,lev=3,rlev=3,ilev=4,lon=4,lon_grd=5,char_dmn_lng80=80,char_dmn_lng26=26,char_dmn_lng04=4,date_dmn=5,fl_dmn=3,lsmlev=6,wvl=2,time_int_udunits=1;time_udunits=3;lon_T42=128,lat_T42=64,lat_times_lon=8,gds_crd=8,gds_ncd=8,lon_cal=10,lat_cal=10,pck_crd=4,vrt_nbr=2,time=10;
// 20231019: Restore NC_UNLIMITED dimension
//dgn=1,bnd=2,lat=2,lat_grd=3,lev=3,rlev=3,ilev=4,lon=4,lon_grd=5,char_dmn_lng80=80,char_dmn_lng26=26,char_dmn_lng04=4,date_dmn=5,fl_dmn=3,lsmlev=6,wvl=2,time_int_udunits=1;time_udunits=3;lon_T42=128,lat_T42=64,lat_times_lon=8,gds_crd=8,gds_ncd=8,lon_cal=10,lat_cal=10,pck_crd=4,vrt_nbr=2,time=unlimited;
// 20231020: Temporarily eliminate NC_UNLIMITED dimension so NCO 5.1.9+ distribution does not break when building with netCDF <= 4.9.2
dgn=1,bnd=2,lat=2,lat_grd=3,lev=3,rlev=3,ilev=4,lon=4,lon_grd=5,char_dmn_lng80=80,char_dmn_lng26=26,char_dmn_lng04=4,date_dmn=5,fl_dmn=3,lsmlev=6,wvl=2,time_int_udunits=1;time_udunits=3;lon_T42=128,lat_T42=64,lat_times_lon=8,gds_crd=8,gds_ncd=8,lon_cal=10,lat_cal=10,pck_crd=4,vrt_nbr=2,time=10;
 variables:
  :Conventions = "CF-1.5";
  :history = "History global attribute.\nTextual attributes like history often have embedded newlines like this.\nSuch newlines should serve as linebreaks on the screen to enhance legibility like this.\nFriendly CDL converters print a single NC_CHAR attribute as a comma-separated list of strings where each embedded delimiter marks a linebreak. This makes poetry embedded in CDL much nicer to read (except for the printed literal \\n\'s---those are an eyesore):\n\nA POET by Hafiz\n\nA poet is someone\nWho can pour light into a cup,\nThen raise it to nourish\nYour beautiful parched, holy mouth\n";
  :lorem_ipsum = "The Lorem Ipsum attribute demonstrates the legibility of text without embedded linebreaks:\nLorem ipsum dolor sit amet, consectetur adipiscing elit, sed do eiusmod tempor incididunt ut labore et dolore magna aliqua. Ut enim ad minim veniam, quis nostrud exercitation ullamco laboris nisi ut aliquip ex ea commodo consequat. Lady Gaga amat indueris vestimento laetus. Duis aute irure dolor in reprehenderit in voluptate velit esse cillum dolore eu fugiat nulla pariatur. Excepteur sint occaecat cupidatat non proident, sunt in culpa qui officia deserunt mollit anim id est laborum.";
  :julian_day = 200000.04;
  :RCS_Header = "$Header$";
  string :sng_att = "Test global string attribute"; // 20130723 This is how to specify global string attributes

//	netCDF4-only atomic types
	int64 int64_var_max;
	int64_var_max:long_name = "int64-type variable";

	int64 int64_var;
	int64_var:long_name = "int64-type variable";

	string string_var;
	string_var:long_name = "string-type variable";

	string string_var2;
	string_var2:long_name = "string-type variable with default XML separator";

	string string_arr_var(lon);
	string_arr_var:long_name = "arrays of string-types";   

	string string_greek(lat,lon);
	string_greek:long_name = "2D arrayof string-types";   

	ubyte ubyte_var;
	ubyte_var:long_name = "ubyte-type variable";

	uint uint_var_max;
	uint_var_max:long_name = "uint-type variable";

	uint uint_var;
	uint_var:long_name = "uint-type variable";

	uint64 uint64_var;
	uint64_var:long_name = "uint64-type variable";

	ushort ushort_var;
	ushort_var:long_name = "ushort-type variable";

//	netCDF3 atomic types:
	int date_int(date_dmn);
	date_int:long_name = "Date (as array of ints: YYYY,MM,DD,HH,MM)";

	float dgn(dgn);
	dgn:long_name = "degenerate coordinate (dgn means degenerate, i.e., of size 1)";

	float dgn_var(dgn);
	dgn_var:long_name = "degenerate variable (dgn means degenerate, i.e., of size 1)";

	float lat(lat);
	lat:long_name = "Latitude (typically midpoints)";
	lat:units = "degrees_north";
	lat:bounds = "lat_bnd";

	float lat_bnd(lat,vrt_nbr);
	lat_bnd:purpose = "Cell boundaries for lat coordinate";

	float lat_grd(lat_grd);
	lat_grd:long_name = "Latitude grid (typically interfaces)";
	lat_grd:units = "degrees_north";

	float lat_cpy(lat);
	float lev_cpy(lev);
	float lat_var(lat);
	float lat_wgt(lat);
	float lon_T42(lon_T42);
	float lat_T42(lat_T42);

	float lat_1D_rct(lat_times_lon);
	lat_1D_rct:long_name = "Latitude for 2D rectangular grid stored as 1D arrays";
	lat_1D_rct:units = "degrees_north";

	float lon_1D_rct(lat_times_lon);
	lon_1D_rct:long_name = "Longitude for 2D rectangular grid stored as 1D arrays";
	lon_1D_rct:units = "degrees_east";

	float lat_1D_rrg(lat_times_lon);
	lat_1D_rrg:long_name = "Latitude for 2D irregular grid stored as 1D arrays";
	lat_1D_rrg:units = "degrees_north";

	float lon_1D_rrg(lat_times_lon);
	lon_1D_rrg:long_name = "Longitude for 2D irregular grid stored as 1D arrays";
	lon_1D_rrg:units = "degrees_east";

	int lat_times_lon(lat_times_lon);
	lat_times_lon:long_name = "Element index (i.e., C-based storage order) for 2D coordinate grids stored as 1D arrays";

        float lat_2D_rct(lat,lon);
	lat_2D_rct:long_name = "Latitude for 2D rectangular grid stored as 2D array";
	lat_2D_rct:units = "degrees_north";

	float lon_2D_rct(lat,lon);
	lon_2D_rct:long_name = "Longitude for 2D rectangular grid stored as 2D array";
	lon_2D_rct:units = "degrees_east";

	float lat_2D_rrg(lat,lon);
	lat_2D_rrg:long_name = "Latitude for 2D irregular grid stored as 2D array";
	lat_2D_rrg:units = "degrees_north";

	float lon_2D_rrg(lat,lon);
	lon_2D_rrg:long_name = "Longitude for 2D irregular grid stored as 2D array";
	lon_2D_rrg:units = "degrees_east";

	int lat_times_lon_nbr;
	lat_times_lon_nbr:long_name = "Number of elements in 2D coordinate grids. Rectangular and irregular test grids have this many total elements. The coordinates and elements are stored as 1D or 2D arrays for grid types 1D and 2D respectively.";

	float lev(lev);
	lev:purpose = "Monotonically increasing coordinate pressure";
	lev:long_name = "hybrid level at midpoints (1000*(A+B))";
	lev:units = "hPa";
	lev:positive = "down";
	lev:A_var = "hyam";
	lev:B_var = "hybm";
	lev:P0_var = "P0";
	lev:PS_var = "PS";
	lev:bounds = "lev_bnd";
        lev:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate";
        lev:formula_terms = "a: hyam b: hybm p0: P0 ps: PS";
        lev:formula_readable = "prs_mdp[time,lat,lon,lev]=P0*hyam+PS*hybm";

	float ilev(ilev);
	ilev:purpose = "Monotonically increasing coordinate pressure";
	ilev:long_name = "hybrid level at interfaces (1000*(A+B))";
	ilev:units = "hPa";
	ilev:positive = "down";
	ilev:A_var = "hyai";
	ilev:B_var = "hybi";
	ilev:P0_var = "P0";
	ilev:PS_var = "PS";
        ilev:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate";
        ilev:formula_terms = "a: hyai b: hybi p0: P0 ps: PS";
        ilev:formula_readable = "prs_ntf[time,lat,lon,ilev]=P0*hyai+PS*hybi";

	float lev_bnd(lev,vrt_nbr);
	lev_bnd:purpose = "Cell boundaries for lev coordinate";

 	float rlev(rlev);
	rlev:purpose = "Monotonically decreasing coordinate pressure";

	float lon(lon);
	lon:long_name = "Longitude (typically midpoints)";
	lon:units = "degrees_east";

	// 20220827: Lat and Lon dimensions break NCZarr->POSIX writes such as
	// ncea -O -C -v lon,three_dmn_rec_var,time,time_bnds,climatology_bounds file:///Users/zender/nco/data/h0001#mode=nczarr,file ~/out.nc
	// Case-insensitive matching of dimension IDs may be at play?
	// Eliminating Lat/Lon dimensions fixes the issue
	//double Lon(Lon);
	double Lon(lon);
	Lon:long_name = "Longitude";
	Lon:units = "degrees";
	Lon:purpose = "Longitude coordinate originally stored as -180 to 180";
	Lon:notes = "Longitude = [-180.0,180.0) is not CF-compliant, yet is common";

	//double LatLon(Lat,Lon);
	double LatLon(lat,lon);
	LatLon:long_name = "2D variable originally stored on -180 to 180 longitude grid";
	LatLon:units = "fraction";
	LatLon:purpose = "Demonstrate remapping of [-180,180) to [0,360) longitude-grid data";

	//double Lat(Lat);
	double Lat(lat);
	Lat:long_name = "Latitude";
	Lat:units = "degrees_north";
	Lat:purpose = "Latitude paired with Longitude coordinate originally stored as -180 to 180.";

	double lond(lon);
	lond:long_name = "Longitude (typically midpoints), double precision";
	lond:units = "degrees_east";

	float lonf(lon);
	lonf:long_name = "Longitude (typically midpoints), single precision";
	lonf:units = "degrees_east";

	float lon_grd(lon_grd);
	lon_grd:long_name = "Longitude grid (typically interfaces)";
	lon_grd:units = "degrees_east";

	double time(time);
	time:long_name = "time";
	time:units = "days since 1964-03-12 12:09:00 -9:00"; 
	time:calendar = "gregorian";
	time:bounds = "time_bnds";
	time:climatology = "climatology_bounds";

	float time_bnds(time,vrt_nbr);
	time_bnds:purpose = "Cell boundaries for time coordinate";

	float climatology_bounds(time,vrt_nbr);
	climatology_bounds:purpose = "Variable containing CF-compliant climatology bounds for time dimension";

	double time_rpt(time);
	time_rpt:long_name = "A repeating sequence to check compliance of MRO";
	time_rpt:purpose = "Sequence is 1,2,3,1,2,3,1,2,3,1. Average of every third element should be the same as the element, e.g., ncra -O --mro -d time,,,3,3 ~/nco/data/in.nc ~/foo.nc;ncks -C -v time_rpt ~/foo.nc";

        double lon_cal(lon_cal);
	lon_cal:long_name = "lon_cal";
	lon_cal:units = "days since 1964-2-28"; 
	lon_cal:calendar = "365_day";

	double lat_cal(lat_cal);
	lat_cal:long_name = "lat_cal";
	lat_cal:units = "days since 1964-2-28"; 
	lat_cal:calendar = "360_day";

	double tm_scn;
        tm_scn:units = "seconds since 2013-01-01";

	double tm_std;
        tm_std:units = "days since 2013-01-01";

	double tm_grg;
        tm_grg:units = "days since 2013-01-01";
        tm_grg:calendar = "gregorian"; // Same as "standard"

	double tm_jln;
        tm_jln:units = "days since 2013-01-01";
        tm_jln:calendar = "julian";

	double tm_360;
        tm_360:units = "days since 2013-01-01";
        tm_360:calendar = "360_day";

	double tm_365;
        tm_365:units = "days since 2013-01-01";
        tm_365:calendar = "365_day"; // Same as "noleap"

	double tm_366;
        tm_366:units = "days since 2013-01-01";
        tm_366:calendar = "366_day"; // Same as "all_leap"

	float lsmlev(lsmlev);
	lsmlev:purpose = "Homebrew level coordinate for LSM";
	lsmlev:long_name = "Soil depth";
	lsmlev:units = "meter";

	float wvl(wvl);
	wvl:long_name = "Wavelength";
	wvl:units = "meter";

	int od(time);

	double areacella(lat,lon);
        areacella:standard_name = "area";
        areacella:long_name = "area";
	areacella:units = "meter2";
	areacella:purpose = "Variable to hold cell areas of 2D fields. Intended to be pointed to by cell_measures attribute of 2D fields. Would have named it plain-old area but too many regression tests already depend on 1D float area below. areacella is name used by ESGF-distributed versions of some CESM simulations anyway, e.g., baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_atmos_fx_CCSM4_amip_r0i0p0.nc areacella: areacella_fx_CCSM4_amip_r0i0p0.nc";

	float area(lat);
	area:long_name = "area";
	area:units = "meter2";

	float area2(lat);
	area2:long_name = "area version 2";
	area2:units = "meter2";

	float area_asm(lat);
	area_asm:long_name = "area asymmetric";
	area_asm:units = "meter2";

	float hyam(lev);
	hyam:long_name = "hybrid A coefficient at layer midpoints";

	float hybm(lev);
	hybm:long_name = "hybrid B coefficient at layer midpoints";

	float hyai(ilev);
	hyai:long_name = "hybrid A coefficient at layer interfaces";

	float hybi(ilev);
	hybi:long_name = "hybrid B coefficient at layer interfaces";

	float P0;
	P0:long_name = "reference pressure";
	P0:units = "pascal";

        float cnv_CF_grd(lat,lon);
	cnv_CF_grd:long_name = "test CF grid_mapping convention";
        cnv_CF_grd:grid_mapping = "albers_conical_equal_area";
        cnv_CF_grd:purpose = "Test whether grid_mapping is propagated with coordinate";

        char mapping;
        mapping:geoid = "eigen-6c4" ;
	mapping:grid_mapping_name = "polar_stereographic" ;
	mapping:latitude_of_projection_origin = -90. ;
	mapping:standard_parallel = -71. ;
	mapping:straight_vertical_longitude_from_pole = 0. ;
	mapping:semi_major_axis = 6378273. ;
	mapping:inverse_flattening = 298.27940504282 ;
	mapping:false_easting = 0. ;
	mapping:false_northing = 0. ;

        char albers_conical_equal_area;
        albers_conical_equal_area:long_name = "Albers Conical Equal Area Projection";
        albers_conical_equal_area:purpose = "Test that this grid_mapping is propagated with all associated variables (like cnv_CF_grd)";
        albers_conical_equal_area:grid_mapping_name = "albers_conical_equal_area";
        albers_conical_equal_area:false_easting = 0.;
        albers_conical_equal_area:false_northing = 0.;
        albers_conical_equal_area:latitude_of_projection_origin = 40.;
        albers_conical_equal_area:longitude_of_central_meridian = -101.;
        albers_conical_equal_area:standard_parallel = 20., 60.;
        albers_conical_equal_area:longitude_of_prime_meridian = 0.;
        albers_conical_equal_area:semi_major_axis = 6378137.;

	float cnv_CF_crd(gds_crd);
	cnv_CF_crd:long_name = "test CF coordinates conventions";
	cnv_CF_crd:coordinates = "lat_gds lon_gds ";
	cnv_CF_crd:reason = "Test whether coordinates attribute strings that end with a space break after nco_var_lst_crd_ass_add() call to nco_lst_prs_2d()";

	float cnv_CF_ncl(time);
	cnv_CF_ncl:long_name = "test CF ancillary_variables convention";
        cnv_CF_ncl:standard_name = "specific_humidity";
        cnv_CF_ncl:ancillary_variables = "cnv_CF_ncl_var_1 cnv_CF_ncl_var_2";
        cnv_CF_ncl:purpose = "Main variable that has ancillary variables named cnv_CF_ncl_var_1 and cnv_CF_ncl_var_2";

	float cnv_CF_ncl_var_1(time);
	cnv_CF_ncl_var_1:long_name = "test CF ancillary_variables convention";
        cnv_CF_ncl_var_1:standard_name = "specific_humidity standard_error";
        cnv_CF_ncl_var_1:purpose = "Ancillary variable for cnv_CF_ncl. Other ancillary variable is cnv_CF_ncl_var_2.";

	float cnv_CF_ncl_var_2(time);
	cnv_CF_ncl_var_2:long_name = "test CF ancillary_variables convention";
        cnv_CF_ncl_var_2:standard_name = "specific_humidity detection_limit";
        cnv_CF_ncl_var_2:purpose = "Ancillary variable for cnv_CF_ncl. Other ancillary variable is cnv_CF_ncl_var_1.";

	float PS(time,lat,lon);
	PS:long_name = "surface pressure";
	PS:units = "pascal";

	char fl_dmn(fl_dmn);
	fl_dmn:long_name = "Character coordinate";
	fl_dmn:units = "[chr]";

	double lat_gds(gds_crd);
	lat_gds:long_name = "Latitude";  
	lat_gds:standard_name = "latitude";
	lat_gds:units="degree";
	lat_gds:purpose = "1-D latitude coordinate referred to by geodesic grid variables";

	double lon_gds(gds_crd);
	lon_gds:long_name = "Longitude";
	lon_gds:standard_name = "longitude";
	lon_gds:units="degree";
	lon_gds:purpose = "1-D longitude coordinate referred to by geodesic grid variables";

	float gds_crd(gds_crd);
	gds_crd:long_name = "Geodesic coordinate";
	gds_crd:units = "degree";
	gds_crd:purpose = "enumerated coordinate like those that might define points in a geodesic grid";
	gds_crd:coordinates = "lat_gds lon_gds";

	float gds_var(gds_crd);
	gds_var:long_name = "Geodesic variable";
	gds_var:units = "meter";
	gds_var:purpose = "Test auxiliary coordinates like those that define geodesic grids";
	gds_var:coordinates = "lat_gds lon_gds";

	float gds_3dvar(time,gds_crd);
	gds_3dvar:long_name = "Geodesic variable";
	gds_3dvar:units = "meter";
	gds_3dvar:coordinates = "lat_gds lon_gds";
	gds_3dvar:purpose = "Test auxiliary coordinates like those that define geodesic grids";

	float gds_var_ncd(gds_ncd);
	gds_var_ncd:long_name = "Geodesic variable on non-coordinate grid";
	gds_var_ncd:units = "meter";
	gds_var_ncd:purpose = "Test auxiliary coordinates like those that define geodesic grids but where underlying dimension is a non-coordinate dimension";
	gds_var_ncd:coordinates = "lat_gds_ncd lon_gds_ncd";

	double lat_gds_ncd(gds_ncd);
	lat_gds_ncd:long_name = "Latitude";  
	lat_gds_ncd:standard_name = "latitude";
	lat_gds_ncd:units="degree";
	lat_gds_ncd:purpose = "1-D latitude coordinate referred to by \"non-coordinate\" (ncd) geodesic grid variables";

	double lon_gds_ncd(gds_ncd);
	lon_gds_ncd:long_name = "Longitude";
	lon_gds_ncd:standard_name = "longitude";
	lon_gds_ncd:units="degree";
	lon_gds_ncd:purpose = "1-D longitude coordinate referred to by \"non-coordinate\" (ncd) geodesic grid variables";

	int nbdate;
	nbdate:long_name = "base date as 6- or 8-digit integer (YYMMDD or YYYYMMDD)";

	int date(time);
	date:long_name = "current date as 6- or 8-digit integer (YYMMDD or YYYYMMDD)";

	float lon_wgt(lon);
	lon_wgt:long_name = "Gaussian weights";
	lon_wgt:purpose = "Gaussian weights which sum to two for n = 4. These weights all have floor of 0.0 so should cause SIGFPE when applied to integer types in weighted average.";

	float ppc_flt_2D(time,lat);
        ppc_flt_2D:long_name = "Precision-Preserving Compression, single precision, two dimensional array, negative values";
        ppc_flt_2D:purpose = "test --ppc switches";
        ppc_flt_2D:original_values="-1.0 -- -20.0";

	double ppc_dbl(time);
        ppc_dbl:long_name = "Precision-Preserving Compression, double precision";
        ppc_dbl:purpose = "test --ppc switches";
        ppc_dbl:original_values="0.0,0.1,0.12,0.123,0.1234,0.12345,0.123456,0.1234567,0.12345678,0.123456789";

	float ppc_flt(time);
        ppc_flt:long_name = "Precision-Preserving Compression, single precision";
        ppc_flt:purpose = "test --ppc switches";
        ppc_flt:original_values="0.0,0.1,0.12,0.123,0.1234,0.12345,0.123456,0.1234567,0.12345678,0.123456789";

	double ppc_big(time);
        ppc_big:long_name = "Precision-Preserving Compression, big numbers";
        ppc_big:purpose = "test --ppc switches";
        ppc_big:original_values="123456789e-10,123456789e-9,123456789e-8,123456789e-7,123456789e-6,123456789e-5,123456789e-4,123456789e-3,123456789e-2,123456789e-1";

	float ppc_btg(time);
	ppc_btg:long_name = "Precision-Preserving Compression, bigger numbers";
        ppc_btg:purpose = "test --ppc switches";
        ppc_btg:original_values="1234567890e20,1234567890e19,1234567890e18,1234567890e17,1234567890e16,1234567890e15,1234567890e14,1234567890e13,1234567890e12,1234567890e11";

	float ppc_btg_scl;
        ppc_btg_scl:long_name = "Precision-Preserving Compression, bigger numbers, scalar";
        ppc_btg_scl:purpose = "test --ppc switches";
        ppc_btg_scl:original_value="1234567890e11";

	double ppc_hgh(time);
        ppc_hgh:long_name = "Precision-Preserving Compression, high precision";
        ppc_hgh:purpose = "test --ppc switches";

	double ppc_hgr(time);
        ppc_hgr:long_name = "Precision-Preserving Compression, higher precision";
        ppc_hgr:purpose = "test --ppc switches";

	float ppc_tst(time);
        ppc_tst:long_name = "Precision-Preserving Compression, single precision tests";
        ppc_tst:purpose = "test --ppq";
        ppc_tst:original_values="0.0,_,0.1234567,-0.1234567,64,-64,123456789e25,123456789e-25,3.1415926535897932384626433832795029,-3.1415926535897932384626433832795029";

	float ppc_dcm(time);
        ppc_dcm:long_name = "Precision-Preserving Compression, decimal tests";
        ppc_dcm:purpose = "test --ppq";
        ppc_dcm:original_values="55,155,255,355,455,555,655,755,855,955";

	float qnt_flt_tst1(dgn);
        qnt_flt_tst1:long_name = "Quantization test, single precision";
        qnt_flt_tst1:original_values="1.1111111";

	double qnt_dbl_tst1(dgn);
        qnt_dbl_tst1:long_name = "Quantization test, double precision";
        qnt_dbl_tst1:original_values="1.111111111111";

	float qnt_flt_tst2(lon_grd);
        qnt_flt_tst2:long_name = "Quantization test, single precision";
        qnt_flt_tst2:original_values="1.11111111, 1.0, 9.99999999, 12345.67, .1234567";

	double qnt_dbl_tst2(lon_grd);
        qnt_dbl_tst2:long_name = "Quantization test, double precision";
        qnt_dbl_tst2:original_values="1.1111111, 1.0, 9.999999999, 1234567890.12345, 123456789012345.0";

	char md5_a;
	md5_a:long_name = "the letter a";
	md5_a:purpose = "String with known MD5 digest"; 
	md5_a:MD5_known_checksum = "0cc175b9c0f1b6a831c399e269772661"; 

	char md5_abc(lev);
	md5_abc:long_name = "the letters abc";
	md5_abc:purpose = "String with known MD5 digest"; 
	md5_abc:MD5_known_checksum = "900150983cd24fb0d6963f7d28e17f72";

	float msk_prt_mss_prt(lon);
	msk_prt_mss_prt:long_name = "partial mask, partial missing value example";
	msk_prt_mss_prt:_FillValue = 1.0e36f;

	float mss_val(lon);
	mss_val:long_name = "partial missing value example";
	mss_val:_FillValue = 1.0e36f;

	float mss_val_scl;
	mss_val_scl:long_name = "scalar missing value";
	mss_val_scl:_FillValue = 1.0e36f;

	float mss_val_scl_sml;
	mss_val_scl_sml:long_name = "scalar missing value";
	mss_val_scl_sml:purpose = "Unlike mss_val_scl, mss_val_scl_sml has a missing value that fits within any packed data type range";
	mss_val_scl_sml:_FillValue = 1.0e4f;

	float mss_val_fst(lon);
	mss_val_fst:long_name = "offset partial missing value example";
	mss_val_fst:_FillValue = -999.0f;

	float fll_val(lon);
	fll_val:long_name = "_FillValue example";
	fll_val:_FillValue = -999.0f;

	float fll_val_mss_val(lon);
	fll_val_mss_val:long_name = "_FillValue example";
	fll_val_mss_val:_FillValue = -999.0f;
	fll_val_mss_val:missing_value = -999.0f;

	float nan_arr(lat);
	nan_arr:long_name = "Intended for array representation of IEEE NaN";
	nan_arr:note = "20120308 Apparently netCDF ncgen chokes on variable names of nan and NaN";
	nan_arr:note2 = "20120330 netCDF ncgen on AIX/bluefire chokes on variable/attribute values of nan";
	nan_arr:note3 = "20120625 netCDF ncgen on netCDF 4.1.1 on apparently chokes on variable/attribute values of nan";
	nan_arr:note4 = "If your NCO build fails because your version of netCDF does not support nan, then cd to the directory that contains the file nco/data/in.cdl and run the command in note5 first and then try to build again";
	nan_arr:note5 = "sed -e 's/nan;/1.0f;/' in.cdl > foo.cdl;ncgen -b -o in.nc foo.cdl";
	nan_arr:note6 = "It is too troublesome to distribute in.cdl with references to NaNs because users always build with old netCDF versions that do not support it. So just comment out nan's for now.";
	//	nan_arr:_FillValue = nan;
		nan_arr:_FillValue = 1.0f;

	float nan_scl;
	nan_scl:long_name = "Intended for scalar representation of IEEE NaN";
	nan_scl:note = "20120308 Apparently netCDF ncgen chokes on variable names of nan and NaN";
	nan_scl:note2 = "20120330 netCDF ncgen on AIX/bluefire chokes on variable/attribute values of nan";
	nan_scl:note3 = "20120625 netCDF ncgen on netCDF 4.1.1 on apparently chokes on variable/attribute values of nan";
	nan_scl:note6 = "It is too troublesome to distribute in.cdl with references to NaNs because users always build with old netCDF versions that do not support it. So just comment out nan's for now.";
	// nan_scl:_FillValue = nan;
        nan_scl:_FillValue = 1.0f;

	float nm_spc;
	nm_spc:long_name = "Variable name with space (invalid)";

	float nm_pnd;
	nm_pnd:long_name = "Variable name with pound symbol (invalid)";

	float no_mss_val(lon);
	no_mss_val:long_name = "no missing value";

	float val_one_mss(lat);
	val_one_mss:long_name = "one regular value, one missing value";
	val_one_mss:_FillValue = 1.0e36f;

	short rec_var_pck_scale_factor_only(time);
	rec_var_pck_scale_factor_only:long_name = "Array packed with scale factor only";
	rec_var_pck_scale_factor_only:note = "Original packed value was 1s..10s with scale_factor = 10.0d no add_offset. Unpacked value should be 10.0 = 10.0d*1s + 0.0d through 100 = 10.0d*1s + 0.0d. Average value should be 55.";
	rec_var_pck_scale_factor_only:scale_factor = 10.0d;

	short pck;
	pck:long_name = "Scalar variable, double, packed as short";
	pck:note = "Original packed value was 1s with scale_factor = 2.0d and add_offset = 1.0d. Unpacked value (netCDF convention) should be 3.0 = 2.0d*1s + 1.0d. Unpacked value (HDF convention) should be 0.0 = 2.0d*(1s-1.0d). NCO algorithms would pack this variable as scale_factor = 0.0d and add_offset = 3.0d.";
	pck:scale_factor = 2.0d;
	pck:add_offset = 1.0d;

	short pck_3;
	pck_3:long_name = "Scalar variable, double, packed as short";
	pck_3:note = "Original packed value was 1s with scale_factor = 2.0d and add_offset = 1.0d. Unpacked value (netCDF convention) should be 3.0 = 2.0d*1s + 1.0d. Unpacked value (HDF convention) should be 0.0 = 2.0d*(1s-1.0d). NCO algorithms would pack this variable as scale_factor = 0.0d and add_offset = 3.0d.";
	pck_3:scale_factor = 2.0d;
	pck_3:add_offset = 1.0d;

	short pck_5;
	pck_5:long_name = "Scalar variable, double, packed as short";
	pck_5:note = "Original packed value was 2s with scale_factor = 2.0d and add_offset = 1.0d. Unpacked value (netCDF convention) should be 5.0 = 2.0d*2s + 1.0d. Unpacked value (HDF convention) should be 2.0 = 2.0d*(2s-1.0d). NCO algorithms would pack this variable as scale_factor = 0.0d and add_offset = 5.0d.";
	pck_5:scale_factor = 2.0d;
	pck_5:add_offset = 1.0d;

	short pck_7;
	pck_7:long_name = "Scalar variable, double, packed as short";
	pck_7:note = "Original packed value was 1s with scale_factor = 4.0d and add_offset = 3.0d. Unpacked value (netCDF convention) should be 7.0 = 4.0d*1s + 3.0d. Unpacked value (HDF convention) should be -8.0 = 4.0d*(1s-3.0d). NCO algorithms would pack this variable as scale_factor = 0.0d and add_offset = 7.0d.";
	pck_7:scale_factor = 4.0d;
	pck_7:add_offset = 3.0d;

	short pck_arr(lon);
	pck_arr:long_name = "Array variable, double, packed as short";
	pck_arr:note = "Packed value is -32767s, 0s, 1s, 32767s, unpacked is same in double";
	pck_arr:scale_factor = 1.0d;
	pck_arr:add_offset = 0.0d;

	short pck_crd(pck_crd);
	pck_crd:long_name = "Coordinate array variable, float, packed as short";
	pck_crd:note = "Packed value is -32767s, 0s, 1s, 32767s, unpacked is factor of 10 different, offset by 73 in float";
	pck_crd:scale_factor = 10.0f;
	pck_crd:add_offset = 73.0f;

	double upk;
	upk:long_name = "Unpacked scalar variable";
	upk:note = "Unpacked value is 3.0d0, upk=unpack(pck)= 2.0d0*1s + 1.0d0 = 3.0d0. Packing this variable should create an NC_SHORT scalar = 0s with packing attribute add_offset=3.0d and either no scale_factor (ncap) or scale_factor = 0.0d (ncpdq).";

	double upk_arr(lon);
	upk_arr:long_name = "Unpacked array";
	upk_arr:note = "Unpacked value is -32767.d, 0.d, 1.d, 32767.d, packed is same in short. Packing algorithm should yield an NC_SHORT array = [] with packing attributes scale_factor=1.0d, add_offset=0.0d";

	float val_eminusten;
	val_eminusten:long_name = "Floating point number with exponent ending in zero to test sng_trm_trl_zro()";
        val_eminusten:att_eminusten = 1.1e-10f;

	int val_one_int;
	val_one_int:long_name = "scalar integer equal to 1";
	val_one_int:_FillValue = -99l;

	int val_one_one_int(lat);
	val_one_one_int:long_name = "1, 1";
	val_one_one_int:_FillValue = -99l;

	short val_max_max_sht(lat);
	val_max_max_sht:long_name = "17000, 17000";
	val_max_max_sht:_FillValue = -99s;

	int val_one_mss_int(lat);
	val_one_mss_int:long_name = "1, mss_val";
	val_one_mss_int:_FillValue = -99l;

	float val_half;
	val_half:long_name = "Scalar with value 0.5";
	val_half:_FillValue = 1.0e36f;

	float val_half_half(lat);
	val_half_half:long_name = "0.5,0.5";
	val_half_half:_FillValue = 1.0e36f;

	float wgt_one(lat);
	wgt_one:long_name = "all values are one";

	float mss_val_all(lon);
	mss_val_all:long_name = "all missing values example";
	mss_val_all:_FillValue = 1.0e36f;

	float scalar_var;
	scalar_var:long_name = "scalar variable";
	scalar_var:units = "fraction";
	scalar_var:_FillValue = 1.0e36f;

	float float_var;
	float_var:long_name = "float";

	double double_var;
	double_var:long_name = "double";

	double double_var2;
	double_var2:long_name = "double";
	double_var2:_FillValue = 1.0e36;

	double pi;
	pi:long_name = "Pi";
	pi:units = "fraction";

	double pi_arr_dbl(lat,lon);
	pi_arr_dbl:long_name = "Pi array double precision";
	pi_arr_dbl:units = "fraction";
	pi_arr_dbl:original_values = "3.1415926535897932384626433832795029";

	float pi_arr_flt(lat,lon);
	pi_arr_flt:long_name = "Pi array single precision";
	pi_arr_flt:units = "fraction";
	pi_arr_flt:original_values = "3.14159265";

	float pi1(time);
	pi1:long_name = "Pi array single precision starting at pi incremented by 1.0e-6 each element";
        pi1:original_values = "3.1415927, 3.1415937, 3.1415946, 3.1415956, 3.1415966, 3.1415977, 3.1415987, 3.1415997, 3.1416006, 3.1416016";
	
	float pi2(time);
	pi2:long_name = "Pi array single precision starting at pi incremented by 1.0e-6 each element";
        pi2:original_values = "3.1415927, 3.1415937, 3.1415946, 3.1415956, 3.1415966, 3.1415977, 3.1415987, 3.1415997, 3.1416006, 3.1416016";
	
	float pi3(time);
	pi3:long_name = "Pi array single precision starting at pi incremented by 1.0e-6 each element";
        pi3:original_values = "3.1415927, 3.1415937, 3.1415946, 3.1415956, 3.1415966, 3.1415977, 3.1415987, 3.1415997, 3.1416006, 3.1416016";
	
	float pi4(time);
	pi4:long_name = "Pi array single precision starting at pi incremented by 1.0e-6 each element";
        pi4:original_values = "3.1415927, 3.1415937, 3.1415946, 3.1415956, 3.1415966, 3.1415977, 3.1415987, 3.1415997, 3.1416006, 3.1416016";
	
	float pi5(time);
	pi5:long_name = "Pi array single precision starting at pi incremented by 1.0e-6 each element";
        pi5:original_values = "3.1415927, 3.1415937, 3.1415946, 3.1415956, 3.1415966, 3.1415977, 3.1415987, 3.1415997, 3.1416006, 3.1416016";
	
	float pi6(time);
        pi6:long_name = "Pi array single precision starting at pi incremented by 1.0e-6 each element";
        pi6:original_values = "3.1415927, 3.1415937, 3.1415946, 3.1415956, 3.1415966, 3.1415977, 3.1415987, 3.1415997, 3.1416006, 3.1416016";
	
	float pi7(time);
	pi7:long_name = "Pi array single precision starting at pi incremented by 1.0e-6 each element";
        pi7:original_values = "3.1415927, 3.1415937, 3.1415946, 3.1415956, 3.1415966, 3.1415977, 3.1415987, 3.1415997, 3.1416006, 3.1416016";
	
	int int_var;
	int_var:long_name = "int";

	// 20210406: netCDF 4.8.0 no longer supports CDL type "long" as synonym for "int"
	// Uncomment next line to demonstrate backwards-incompatibility of 4.8.0
	//long long_var;
	int long_var;
	long_var:long_name = "long";
	long_var:purpose = "Variable of CDL type=long, which is deprecated for int. Included to test back-compatibility";
	long_var:notes = "This check will fail with netCDF 4.8.0 if CDL type of variable is long not int. This failure with 4.8.0 was fixed in netCDF master within a few weeks and the problem should not be present in subsequent  (or prior) netCDF versions.";

	short short_var;
	short_var:long_name = "short";

	char char_var;
	char_var:long_name = "char";

	char char_var_space;
	char_var_space:long_name = "Character variable with whitespace on ends";

	char char_var_nul;
	char_var_nul:long_name = "Character variable containing one NUL specified as empty string: \"\"";

	char char_var_nul_c_format;
	char_var_nul_c_format:long_name = "Character variable containing one NUL specified in C-format: \'\\0\'";

	char char_var_zero;
	char_var_zero:long_name = "Character variable containing zero";

	char char_var_1D_arr(time);
        char_var_1D_arr:long_name = "char-type 1D variable array";

	char char_var_2D_arr(lat,lon);
        char_var_2D_arr:long_name = "char-type 2D variable array";
	
        // 20131015: This confuses the XML parser. Omit it for now.
	// char char_var_multinul(lev);
	// char_var_multinul:long_name = "Character variable containing multiple NULs";

	char fl_nm(char_dmn_lng80);
	fl_nm:long_name = "Variable contains a file name";

	char fl_nm_arr(fl_dmn,char_dmn_lng80);
	fl_nm_arr:long_name = "Variable that contains a short array of file names";
	fl_nm_arr:units = "[sng]";

	char fl_nm_rec(time,char_dmn_lng80);
	fl_nm_rec:long_name = "A record variable of file names";
	fl_nm_rec:units = "[sng]";

	char date_sng(char_dmn_lng26);
	date_sng:long_name = "A single date string";
	date_sng:units = "[sng]";

	char date_rec(time,char_dmn_lng26);
	date_rec:long_name = "A record variable of date strings";
	date_rec:units = "[sng]";

	char non_nul_trm_char_one_dmn(char_dmn_lng04);
	non_nul_trm_char_one_dmn:long_name = "Variable contains a one-dimensional array of characters that is not NUL-terminated";
	non_nul_trm_char_one_dmn:units = "[chr]";

	char non_nul_trm_char_two_dmn(fl_dmn,char_dmn_lng04);
	non_nul_trm_char_two_dmn:long_name = "Variable contains a two-dimensional array of characters that are not NUL-terminated";
	non_nul_trm_char_two_dmn:units = "[chr]";

	byte byt_arr(lat,lon);
	byt_arr:long_name = "byte array";

	byte byt_2D(lat,lon);

	byte byt_3D(lat,lev,lon);

	byte byt_3D_rec(time,lat,lon);

	byte byt_bln_3D_rec(time,lat,lon);

	byte byte_var;
	byte_var:long_name = "byte";

	byte byte_var_neg;
	byte_var_neg:long_name = "negative byte";

	float zero;
	zero:long_name = "zero";

	float ppc_zro_flt(time);
	ppc_zro_flt:long_name = "array of single precision floating point zeros";

	double ppc_zro_dbl(time);
	ppc_zro_dbl:long_name = "array of double precision floating point zeros";

	int ppc_zro_int(time);
	ppc_zro_int:long_name = "array of integer zeros";

	float one;
	one:long_name = "one";

	float two;
	two:long_name = "two";

	double e_dbl;
	e_dbl:long_name = "e, natural logarithm base";

	float e_flt;
	e_flt:long_name = "e, natural logarithm base";

	float three;
	three:long_name = "three";

	float four;
	four:long_name = "four";

	float negative_one;
	negative_one:long_name = "negative one";

	float lev_var(lev);
	lev_var:long_name = "lev_var";

	float lev_wgt(lev);
	lev_wgt:long_name = "lev_wgt";

	float g;
	g:long_name = "g";

	float grv_sfc;
	grv_sfc:long_name = "Surface gravity on Earth";
	grv_sfc:units = "meter second-2";

	float vmr_CO2;
	vmr_CO2:long_name = "Volumetric mixing ratio of CO2";
	vmr_CO2:units = "molecule molecule-1";

	float mmr_CO2;
	mmr_CO2:long_name = "Mass mixing ratio of CO2";
	mmr_CO2:units = "kilogram kilogram-1";

	float dps_dry;
	dps_dry:long_name = "Dry Deposition";

	float dps_wet;
	dps_wet:long_name = "Wet Deposition";

	float dps_ttl;
	dps_ttl:long_name = "Total Deposition";

	float z(lev);
	z:long_name = "Height";
	z:units = "meter";
	z:purpose = "Height stored with a monotonically increasing coordinate";

	float rz(rlev);
	rz:long_name = "Height";
	rz:units = "meter";
	rz:purpose = "Height stored with a monotonically decreasing coordinate";

	float one_dmn_var(bnd);

	int one_dmn_int_val_one(lat);
	int one_dmn_int_val_two(lat);

	float att_var(time);
	att_var:byte_att = '\000','\001','\002','\177','\200','\201','\376','\377';
	att_var:char_att = "Sentence one.\nSentence two.\n";
	att_var:char_att2 = "Character string containing default XML separator: *|*\n";
	att_var:short_att = 37s;
	att_var:int_att = 73;
        att_var:float_att = 73.0f,72.0f,71.0f,70.010f,69.0010f,68.010000f,67.01000100f;
	att_var:double_att = 73.0,72.0,71.0,70.010,69.0010,68.010000,67.01000100;
	att_var:ubyte_att = 0ub, 1ub, 2ub, 127ub, 128ub, 254ub, 255ub, 0ub; // 20130712: ncgen 4.3.0 translates this to byte
        att_var:ushort_att = 37us;
        att_var:uint_att = 73ul; // 20161110: ncgen requires "ul" for uint (a simple "u" is interpretd as uint64)
	att_var:int64_att = 9223372036854775807ll; // 20130712: ncgen 4.3.0--4.3.3.1 choke on ll, LL suffix for int64 attributes, and translates -l suffixed numbers to NC_UINT64. Bug reported (netCDF #HEX-795132) and fixed in snapshot 20131117
        att_var:uint64_att = 18446744073709551615ull; // 20130712: ncgen 4.3.0--4.3.3.1 chokes on ull, ULL suffix for uint64 attributes. 20131120: XML treats unsigned as signed types, so toolsui produces errors when reading maximum uint64 values (though not when reading maximum ubyte, ushort, and uint values)
	att_var:string_att1 = "20130723: ncgen -k netCDF-4 version 4.0.x converts quoted string to NC_STRING not NC_CHAR. Incompatible with classic behavior.";
	att_var:string_att2 = "20130712: ncgen -k netCDF-4 version 4.2.x+ converts quoted string to NC_CHAR not NC_STRING. Backwards compatible with classic behavior.";
	string att_var:string_att3 = "20130723: Prefixing full attribute name with \"string\" causes CDL to produce NC_STRING.";
	string att_var:string_att4 = "20130723: Arrays of NC_STRING are simply separated by commas.","If there are commas within a string, well, then, be careful. Did we \"jump the shark\"?","This array comprises three elements. Each is a sentence or three long.";
	string att_var:string_att5 = "20131121: This NC_STRING contains NCO's default XML string separator, *. And it contains multiple sequential copies of that separator, ***. Be sure ncks automatically switches to a different separator, aka the backup separator, the string obtained by removing the two spaces from this:\"* | *\".";

	int att_var_jsn;
        // 20210512: HDF4 ncgen fails on character attributes with whitespace
	att_var_jsn:char\ att\ with\ whitespace = "cf-json.org <http://cf-json.org>";
        att_var_jsn:double\ att\ with\ whitespace = 3.14;
        att_var_jsn:int\ att\ with\ whitespace = 1;
        att_var_jsn:int_array\ att\ with\ whitespace = 1,2;

	// Purpose: Test special characters in names
	// Most special characters need backslash protection
	int att_var_spc_chr;
	att_var_spc_chr:space\ in\ name = "foo";
	att_var_spc_chr:comma_in_name\, = "foo";
	att_var_spc_chr:lt_in_name\< = "foo";
	att_var_spc_chr:gt_in_name\> = "foo";
	att_var_spc_chr:hash_in_name\# = "foo";
	att_var_spc_chr:xclaim_in_name\! = "foo";
	att_var_spc_chr:dollar_in_name\$ = "foo";
	att_var_spc_chr:ampersand_in_name\& = "foo";
	att_var_spc_chr:equals_in_name\= = "foo";
	att_var_spc_chr:semicolon_in_name\; = "foo";
	att_var_spc_chr:colon_in_name\: = "foo";
	att_var_spc_chr:lbrace_in_name\{ = "foo";
	att_var_spc_chr:rbrace_in_name\} = "foo";
	att_var_spc_chr:lparen_in_name\( = "foo";
	att_var_spc_chr:rparen_in_name\) = "foo";
	att_var_spc_chr:lbracket_in_name\[ = "foo";
	att_var_spc_chr:rbracket_in_name\] = "foo";
	att_var_spc_chr:plus_in_name+ = "foo";
	//  : period_in_name. = "foo"; // Likely to cause DAP server error
	att_var_spc_chr:hyphen_in_name- = "foo";
	att_var_spc_chr:at_in_name@ = "foo";

	// Purpose test special chars in char atts 
        int att_sng;
        att_sng:nul_sng = '\0';
	att_sng:empty_sng = "";
        att_sng:space_sng = " ";
	att_sng:zero_sng = "0";
	
	int bnd_var(lev,bnd);
	bnd_var:byte_att = '\0';
	bnd_var:char_att = "Sentence one.\nSentence two.\n";
	bnd_var:short_att = 37s;
	bnd_var:int_att = 73;
	bnd_var:long_att = 73;
	bnd_var:float_att = 73.f;
	bnd_var:double_att = 73.d;

	float three_dmn_var(lat,lev,lon);
	three_dmn_var:long_name = "three dimensional variable with CCM coordinate convention C=[lat,lev,lon], Fortran=(lon,lev,lat)";
	three_dmn_var:units = "fraction";

	float three_dmn_var_crd(lev,lat,lon);
	three_dmn_var_crd:long_name = "three dimensional variable with COORDS coordinate convention C=[lev,lat,lon], Fortran=(lon,lat,lev)";
	three_dmn_var_crd:units = "fraction";

	float three_dmn_var_cf(lev,lat,lon);
	three_dmn_var_cf:long_name = "three dimensional variable with CF \"coordinates\" convention";
	three_dmn_var_cf:coordinates = "lat lev lon";
	three_dmn_var_cf:units = "fraction";

	float three_dmn_var_cf2(lev,lat,lon);
	three_dmn_var_cf2:long_name = "three dimensional variable with CF \"coordinates\" convention for wrong coordinates";
	three_dmn_var_cf2:coordinates = "x y z";
	three_dmn_var_cf2:units = "fraction";

	float prs_sfc(time,lat,lon);
	prs_sfc:long_name = "Surface pressure";
	prs_sfc:units = "pascal";

	float H2O;
	float H2OH2O;
	float H2SO4;
	float H2O_lqd;
	float H2O_ice;
	float Q;
	float Q1;
	float AQ01;
	float QQ01;
	float QA01;
	float Q01Q;
	float Q01;
	float Q02;
	float Q03;
	float Q04;
	float Q05;
	float Q06;
	float Q07;
	float Q08;
	float Q09;
	float Q10;
	float Q11;
	float Q12;
	float Q13;
	float Q14;
	float Q15;
	float Q16;
	float Q17;
	float Q18;
	float Q19;
	float Q20;
	float Q21;
	float Q22;
	float Q23;
	float Q24;
	float Q25;
	float Q26;
	float Q27;
	float Q28;
	float Q29;
	float Q30;
	float Q31;
	float Q32;
	float Q33;
	float Q34;
	float Q35;
	float Q36;
	float Q37;
	float Q38;
	float Q39;
	float Q40;
	float Q41;
	float Q42;
	float Q43;
	float Q44;
	float Q45;
	float Q46;
	float Q47;
	float Q48;
	float Q49;
	float Q50;
	float Q51;
	float Q52;
	float Q53;
	float Q54;
	float Q55;
	float Q56;
	float Q57;
	float Q58;
	float Q59;
	float Q60;
	float Q61;
	float Q62;
	float Q63;
	float Q64;
	float Q65;
	float Q66;
	float Q67;
	float Q68;
	float Q69;
	float Q70;
	float Q71;
	float Q72;
	float Q73;
	float Q74;
	float Q75;
	float Q76;
	float Q77;
	float Q78;
	float Q79;
	float Q80;
	float Q81;
	float Q82;
	float Q83;
	float Q84;
	float Q85;
	float Q86;
	float Q87;
	float Q88;
	float Q89;
	float Q90;
	float Q91;
	float Q92;
	float Q93;
	float Q94;
	float Q95;
	float Q96;
	float Q97;
	float Q98;
	float Q99;
	float Q100;

	float two_dmn_var(lat,lev);
	two_dmn_var:long_name = "two dimensional variable";
	two_dmn_var:units = "fraction";

	float var_msk(lat,lon);
	var_msk:long_name = "Float field for testing masks and wheres";
	var_msk:units = "fraction";

	float var_mss_nil(lon);
        var_mss_nil:purpose = "Test mismatched missing values in variables, masks, and weights. Missing no elements.";
	var_mss_nil:_FillValue = 1.0e36f;

	float var_mss_0(lon);
        var_mss_0:purpose = "Test mismatched missing values in variables, masks, and weights. Missing element index 0.";
	var_mss_0:_FillValue = 1.0e36f;

	float var_mss_1(lon);
        var_mss_1:purpose = "Test mismatched missing values in variables, masks, and weights. Missing element index 1.";
	var_mss_1:_FillValue = 1.0e36f;

	float var_mss_2(lon);
        var_mss_2:purpose = "Test mismatched missing values in variables, masks, and weights. Missing element index 2.";
	var_mss_2:_FillValue = 1.0e36f;
	
	float var_mss_3(lon);
        var_mss_3:purpose = "Test mismatched missing values in variables, masks, and weights. Missing element index 3.";
	var_mss_3:_FillValue = 1.0e36f;
	
	float mask(lat,lon);
	mask:long_name = "Purpose is to mask a variable like ORO";
	mask:units = "fraction";

	float ORO(lat,lon);
	ORO:long_name = "Orography, an enumerated yet continuous type: ocean=0.0, land=1.0, sea ice=2.0";
	ORO:units = "fraction";

	float orog(lat,lon);
	orog:long_name = "Orography, an enumerated yet continuous type: ocean=0.0, land=1.0, sea ice=2.0";
	orog:units = "fraction";
        orog:original_name = "ORO" ;
        orog:cell_measures = "area: areacella" ;
        orog:purpose = "Replicate processing of files produced by CESM and distributed on ESGF" ;

	float orog2(lat,lon);
	orog2:long_name = "Value of 1 everywhere on latxlon grid";
	orog2:units = "fraction";
        orog2:purpose = "debug TODO nco1138" ;

	float orog3(lat,lon);
	orog3:long_name = "Value of 0 first half, 1 second half on latxlon grid";
	orog3:units = "fraction";
        orog3:purpose = "debug TODO nco1138" ;

	float weight(lat);
	weight:long_name = "Gaussian weight";
	weight:units = "fraction";

	float gw(lat);
	gw:long_name = "gw variable like gw";
	gw:units = "fraction";

	float gw_T42(lat_T42);
	gw_T42:long_name = "gw variable like gw_T42";
	gw_T42:units = "fraction";

	float rec_var_flt(time);
	rec_var_flt:long_name = "record variable, float";

	double rec_var_dbl(time);
	rec_var_dbl:long_name = "record variable, double";

	int one_dmn_rec_var(time);
	one_dmn_rec_var:long_name = "one dimensional record variable";
	one_dmn_rec_var:coordinates = "time";
	one_dmn_rec_var:units = "kelvin";

	double one_dmn_rec_wgt(time);
	one_dmn_rec_wgt:long_name = "one dimensional record variable weight";
	
	int one_dmn_rec_var_mdn(time);
	one_dmn_rec_var_mdn:long_name = "one dimensional record variable to test median";
        
	int one_dmn_rec_var_mdn__FillValue(time);
	one_dmn_rec_var_mdn__FillValue:long_name = "one dimensional record variable to test median with _FillValue";
	one_dmn_rec_var_mdn__FillValue:_FillValue = -999;
        
	int one_dmn_rec_var_unsorted(time);
	one_dmn_rec_var_unsorted:long_name = "one dimensional record variable, unsorted";
        
	float one_dmn_rec_var_flt(time);
	one_dmn_rec_var_flt:long_name = "one dimensional record variable, single precision";
        
	float one_dmn_rec_var_flt_mss(time);
	one_dmn_rec_var_flt_mss:long_name = "one dimensional record variable, single precision, missing values";
	one_dmn_rec_var_flt_mss:_FillValue = 1.0e36f;
        
	float one_dmn_rec_var_flt_scl(time);
	one_dmn_rec_var_flt_scl:long_name = "one dimensional record variable, single precision, scaled";
	one_dmn_rec_var_flt_scl:scale_factor = 1.0f;
        
	float one_dmn_rec_var_flt_mss_scl(time);
	one_dmn_rec_var_flt_mss_scl:long_name = "one dimensional record variable, single precision, missing values, scaled";
	one_dmn_rec_var_flt_mss_scl:scale_factor = 1.0f;
	one_dmn_rec_var_flt_mss_scl:_FillValue = 1.0e36f;
        
	float one_dmn_rec_var_dbl(time);
	one_dmn_rec_var_dbl:long_name = "one dimensional record variable, double precision";
	one_dmn_rec_var_dbl:units = "second";
        
	float one_dmn_rec_var_missing_value(time);
	one_dmn_rec_var_missing_value:long_name = "One dimensional record variable with missing data indicated by missing_value attribute only. No _FillValue attribute exists.";
	one_dmn_rec_var_missing_value:missing_value = 1.0e36f;

	float one_dmn_rec_var_mss_val(time);
	one_dmn_rec_var_mss_val:long_name = "One dimensional record variable with all missing data.";
	one_dmn_rec_var_mss_val:_FillValue = 1.0e36f;

	float one_dmn_rec_var__FillValue(time);
	one_dmn_rec_var__FillValue:long_name = "One dimensional record variable with missing data indicated by _FillValue attribute only. No missing_value attribute exists.";
	one_dmn_rec_var__FillValue:_FillValue = 1.0e36f;

	float one_dmn_rec_var_unsorted__FillValue(time);
	one_dmn_rec_var_unsorted__FillValue:long_name = "Unsorted, one dimensional record variable with missing data indicated by _FillValue attribute only. No missing_value attribute exists.";
	one_dmn_rec_var_unsorted__FillValue:_FillValue = 1.0e36f;

	float one_dmn_rec_var_mss_val_arr(time);
	one_dmn_rec_var_mss_val_arr:long_name = "One dimensional record variable with missing data indicated by a _FillValue attribute that is an array. This can be tested with ncrcat. 20120905: ncgen chokes on _FillValue arrays and produces this error: _FillValue: must be a single (possibly compound) value. Deprecate the array for normal use since it prevents ncgen from completing. Uncommment following line when testing for compatibility with software changes.";
//	one_dmn_rec_var_mss_val_arr:_FillValue = 1.0f,2.0f,3.0f;
	one_dmn_rec_var_mss_val_arr:_FillValue = 1.0f;

	int RDM(time);
        
	float tpt(time);
	tpt:long_name = "Temperature";
	tpt:units = "kelvin";
	tpt:hieght = "Leave hieght mispelled for NCO User's guide example";

	double tpt_dbl(time);
	tpt_dbl:long_name = "Temperature stored as double precision floating point";
	tpt_dbl:units = "kelvin";

	float tpt_flt(time);
	tpt_flt:long_name = "Temperature stored as single precision floating point";
	tpt_flt:units = "kelvin";

	double rec_var_dbl_mss_val_dbl_upk(time);
	rec_var_dbl_mss_val_dbl_upk:long_name = "record variable, double, with double missing values";
	rec_var_dbl_mss_val_dbl_upk:purpose = "This variable is used to generate the packed variable rec_var_dbl_mss_val_dbl_pck, so its _FillValue should not be out of range, i.e., it should be representable by a short. However, the _FillValue should itself be the same type as the unpacked variable, NC_DOUBLE in this case.";
	rec_var_dbl_mss_val_dbl_upk:_FillValue = -999.;
	rec_var_dbl_mss_val_dbl_upk:missing_value = -999.;

	double rec_var_dbl_mss_val_sht_upk(time);
	rec_var_dbl_mss_val_sht_upk:long_name = "record variable, double, with double missing values";
	rec_var_dbl_mss_val_sht_upk:purpose = "This variable is used to generate the packed variable rec_var_dbl_mss_val_sht_pck, so its _FillValue should not be out of range, i.e., it should be representable by a short. However, the _FillValue should itself be the same type as the unpacked variable, NC_DOUBLE in this case.";
//	Using intended _FillValue type breaks ncgen (with "_FillValue type mismatch")in netCDF 4.1.1 so comment-out for simplicity
//	rec_var_dbl_mss_val_sht_upk:_FillValue = -999s;
	rec_var_dbl_mss_val_sht_upk:_FillValue = -999.0;
	rec_var_dbl_mss_val_sht_upk:missing_value = -999s;

	short rec_var_dbl_mss_val_dbl_pck(time);
	rec_var_dbl_mss_val_dbl_pck:long_name = "record variable, double, packed as short, with double missing values";
	rec_var_dbl_mss_val_dbl_pck:purpose = "Packed version of rec_var_dbl_mss_val_dbl_upk";
//	Using intended _FillValue type breaks ncgen (with "_FillValue type mismatch")in netCDF 4.1.1 so comment-out for simplicity
//	rec_var_dbl_mss_val_dbl_pck:_FillValue = -999.;
	rec_var_dbl_mss_val_dbl_pck:_FillValue = -999s;
	rec_var_dbl_mss_val_dbl_pck:missing_value = -999.;
        rec_var_dbl_mss_val_dbl_pck:scale_factor = -9.15541313801785e-05;
        rec_var_dbl_mss_val_dbl_pck:add_offset = 5.;

	short rec_var_dbl_mss_val_sht_pck(time);
	rec_var_dbl_mss_val_sht_pck:long_name = "record variable, double, packed as short, with short missing values";
	rec_var_dbl_mss_val_sht_pck:purpose = "Packed version of rec_var_dbl_mss_val_sht_upk";
	rec_var_dbl_mss_val_sht_pck:_FillValue = -999s;
	rec_var_dbl_mss_val_sht_pck:missing_value = -999s;
        rec_var_dbl_mss_val_sht_pck:scale_factor = -9.15541313801785e-05;
        rec_var_dbl_mss_val_sht_pck:add_offset = 5.;

	short scl_dbl_pck;
	scl_dbl_pck:long_name = "scalar variable, double, packed";
	scl_dbl_pck:purpose = "Packed version of number with ncdiff subtraction bug";
        scl_dbl_pck:scale_factor = -9.15541313801785e-05;
        scl_dbl_pck:add_offset = 5.;

	float rec_var_flt_mss_val_flt(time);
	rec_var_flt_mss_val_flt:long_name = "record variable, float, with float missing values";
	rec_var_flt_mss_val_flt:_FillValue = 1.0e36f;

	float rec_var_flt_mss_val_flt_all(time);
	rec_var_flt_mss_val_flt_all:long_name = "record variable, float, with float missing values in every position";
	rec_var_flt_mss_val_flt_all:_FillValue = 1.0e36f;

	float rec_var_flt_mss_val_flt_all_but_one(time);
	rec_var_flt_mss_val_flt_all_but_one:long_name = "record variable, float, with float missing values in every position but one";
	rec_var_flt_mss_val_flt_all_but_one:_FillValue = 1.0e36f;

	float rec_var_flt_mss_val_flt_all_but_two(time);
	rec_var_flt_mss_val_flt_all_but_two:long_name = "record variable, float, with float missing values in every position but two";
	rec_var_flt_mss_val_flt_all_but_two:_FillValue = 1.0e36f;

	short rec_var_flt_pck(time);
	rec_var_flt_pck:long_name = "record variable, float, packed into short";
        rec_var_flt_pck:purpose = "Demonstrate that rounding of means of packed data are handled correctly";
        rec_var_flt_pck:scale_factor = 0.1f;
        rec_var_flt_pck:add_offset = 100.0f;

	short rec_var_dbl_pck(time);
	rec_var_dbl_pck:long_name = "record variable, double, packed into short";
        rec_var_dbl_pck:purpose = "Demonstrate that rounding of means of packed data are handled correctly";
        rec_var_dbl_pck:scale_factor = 0.1;
	rec_var_dbl_pck:add_offset = 100.0;
	
	short non_rec_var_flt_pck(lon);
	non_rec_var_flt_pck:long_name = "regular variable, float, packed into short";
        non_rec_var_flt_pck:purpose = "Demonstrate that non-rec dim packed vars are handled correctly";
        non_rec_var_flt_pck:scale_factor = 0.1f;
        non_rec_var_flt_pck:add_offset = 100.0f;

	float rec_var_flt_mss_val_dbl(time);
	rec_var_flt_mss_val_dbl:long_name = "record variable, float, with double missing values";
	rec_var_flt_mss_val_dbl:_FillValue = 1.0e36f;
	rec_var_flt_mss_val_dbl:missing_value = 1.0e36f;
	rec_var_flt_mss_val_dbl:note = "The correct average of this variable is 5.0. The correct sum of this variable is 35.";

	float rec_var_flt_mss_val_int(time);
	rec_var_flt_mss_val_int:long_name = "record variable, float, with integer missing values";
//	Using intended _FillValue type breaks ncgen (with "_FillValue type mismatch")in netCDF 4.1.1 so comment-out for simplicity
//	rec_var_flt_mss_val_int:_FillValue = -999;
	rec_var_flt_mss_val_int:_FillValue = -999.0f;
	rec_var_flt_mss_val_int:missing_value = -999;

	int rec_var_int_mss_val_int(time);
	rec_var_int_mss_val_int:long_name = "record variable, integer, with integer missing values";
	rec_var_int_mss_val_int:_FillValue = -999;

	int rec_var_int_mss_val_flt(time);
	rec_var_int_mss_val_flt:long_name = "record variable, integer, with float missing values";
//	Using intended _FillValue type breaks ncgen (with "_FillValue type mismatch")in netCDF 4.1.1 so comment-out for simplicity
//	rec_var_int_mss_val_flt:_FillValue = -999.0f;
	rec_var_int_mss_val_flt:_FillValue = -999;
	rec_var_int_mss_val_flt:missing_value = -999.0f;

	int rec_var_int_mss_val_dbl(time);
	rec_var_int_mss_val_dbl:long_name = "record variable, integer, with double missing values";
//	Using intended _FillValue type breaks ncgen (with "_FillValue type mismatch")in netCDF 4.1.1 so comment-out for simplicity
//	rec_var_int_mss_val_dbl:_FillValue = -999.0;
	rec_var_int_mss_val_dbl:_FillValue = -999;
	rec_var_int_mss_val_dbl:missing_value = -999.0;

	int rec_var_dbl_mss_val_dbl_pck_lng(time);
	rec_var_dbl_mss_val_dbl_pck_lng:long_name = "record variable, double packed as long, with double missing values";
	rec_var_dbl_mss_val_dbl_pck_lng:purpose = "although not usual, packing doubles into longs (rather than shorts) offers considerable space savings";
//	Using intended _FillValue type breaks ncgen (with "_FillValue type mismatch")in netCDF 4.1.1 so comment-out for simplicity
//	rec_var_dbl_mss_val_dbl_pck_lng:_FillValue = -999.0;
	rec_var_dbl_mss_val_dbl_pck_lng:_FillValue = -999;
	rec_var_dbl_mss_val_dbl_pck_lng:missing_value = -999.0;
        rec_var_dbl_mss_val_dbl_pck_lng:scale_factor = -9.15541313801785e-05;
        rec_var_dbl_mss_val_dbl_pck_lng:add_offset = 5.;

	short rec_var_dbl_mss_val_sht_pck_sht(time);
	rec_var_dbl_mss_val_sht_pck_sht:long_name = "record variable, double packed as short, with short missing values";
	rec_var_dbl_mss_val_sht_pck_sht:_FillValue = -999s;
        rec_var_dbl_mss_val_sht_pck_sht:scale_factor = -9.15541313801785e-05;
	rec_var_dbl_mss_val_sht_pck_sht:add_offset = 5.;

	float rec_var_flt_mss_val_flt_pck_flt(time);
	rec_var_flt_mss_val_flt_pck_flt:long_name = "record variable, float packed as float, with float missing values";
	rec_var_flt_mss_val_flt_pck_flt:purpose = "CESM POP2 ocean model packs SALT, WVEL etc this way";
	rec_var_flt_mss_val_flt_pck_flt:_FillValue = -9.96921e+33;
        rec_var_flt_mss_val_flt_pck_flt:scale_factor = 1000.0;

	float SALT(time);
	SALT:long_name = "record variable, float packed as float, with float missing values";
	SALT:purpose = "CESM POP2 ocean model packs SALT, WVEL etc this way";
	SALT:_FillValue = -9.96921e+33;
        SALT:scale_factor = 1000.0;
	
	char one_dmn_rec_var_sng(time);
	one_dmn_rec_var_sng:long_name = "one dimensional record variable of string";
        one_dmn_rec_var_sng:NB = "20131222: HDF4 ncgen fails on this variable: /usr/bin/hncgen -b -o ~/in.hdf ~/nco/data/in.cdl produces error message that \"string won't fit in this variable\"";

	float time_lon(time,lon);
	time_lon:long_name = "Record variable of longitude coordinate";

	char two_dmn_rec_var_sng(time,lev);
	two_dmn_rec_var_sng:long_name = "two dimensional record variable of string";

	float two_dmn_rec_var(time,lev);
	two_dmn_rec_var:long_name = "two dimensional record variable";
	two_dmn_rec_var:units = "watt meter-2";

	double three_dmn_var_dbl(time,lat,lon);
	three_dmn_var_dbl:long_name = "three dimensional record variable of type double";
	three_dmn_var_dbl:units = "watt meter-2";
	three_dmn_var_dbl:_FillValue = -99.;

	float zg(time,lev,lon);
	zg:long_name = "three dimensional record variable to demonstrate hyperslab bug";
	zg:units = "watt meter-2";
	zg:_FillValue = -99.;

	float three_dmn_rec_var(time,lat,lon);
	three_dmn_rec_var:long_name = "three dimensional record variable";
	three_dmn_rec_var:units = "watt meter-2";
	three_dmn_rec_var:_FillValue = -99.;

	short three_dmn_rec_var_pck(time,lat,lon);
	three_dmn_rec_var_pck:long_name = "three dimensional record variable";
	three_dmn_rec_var_pck:purpose = "should unpack into identical values with three_dmn_rec_var (i.e., 1..80)";
	three_dmn_rec_var_pck:units = "watt meter-2";
	three_dmn_rec_var_pck:_FillValue = -99.;
        three_dmn_rec_var_pck:add_offset = 40.5f ;
        three_dmn_rec_var_pck:scale_factor = -0.001205518f ;

	int three_dmn_var_int(time,lat,lon);
	three_dmn_var_int:long_name = "three dimensional record variable of type int";
	three_dmn_var_int:units = "watt meter-2";
	three_dmn_var_int:_FillValue = -99;
	
	short three_dmn_var_sht(time,lat,lon);
	three_dmn_var_sht:long_name = "three dimensional record variable";
	three_dmn_var_sht:units = "watt meter-2";
	three_dmn_var_sht:_FillValue = -99s;

	int th(time,lat,lon);
	th:long_name = "three dimensional record variable";
	th:units = "watt meter-2";
	th:_FillValue = -99;

	float td(time,dgn);
	td:long_name = "two dimensional record variable stored in td (time,dgn) order (dgn means degenerate, i.e., of size 1)";

	float tx(time,lon);
	tx:long_name = "two dimensional record variable stored in tx (time,lon) order";

	float ty(time,lat);
	ty:long_name = "two dimensional record variable stored in ty (time,lat) order";

	float tz(time,lev);
	tz:long_name = "two dimensional record variable stored in tz (time,lev) order";

	float txyz(time,lon,lat,lev);
	txyz:long_name = "four dimensional record variable stored in txyz (time,lon,lat,lev) order";

	float xyz(lon,lat,lev);
	xyz:long_name = "three dimensional variable stored in xyz (lon,lat,lev) order";
	
	float tyz(time,lat,lev);
	tyz:long_name = "three dimensional record variable stored in tyz (time,lat,lev) order";
	
	float four_dmn_rec_var(time,lat,lev,lon);
	four_dmn_rec_var:long_name = "four dimensional record variable";
	four_dmn_rec_var:units = "watt meter-2";
	four_dmn_rec_var:coordinates = "time lat lev lon";

//	double three_double_dmn(time,lon,lon);
	
	double time_udunits(time_udunits);
	time_udunits:units = "hours since 1900-01-01 00:00:0.0";
	time_udunits:delta_t = "0000-00-00 06:00:0.0";
	time_udunits:purpose = "The dates specified in this variable are ~1999-12-08";

	int time_int_udunits(time_int_udunits);
	time_int_udunits:units = "seconds since 2019-03-12 00:00:00 UTC";
	time_int_udunits:purpose = "time coordinate with integer values to test rebasing";

	float u(time);
	u:long_name = "Zonal wind speed";
	u:units = "meter second-1";

	float v(time);
	v:long_name = "Meridional wind speed";
	v:units = "meter second-1";

	float var_1D_rct(lat_times_lon);
	var_1D_rct:long_name = "Variable for 2D rectangular grid stored as 1D arrays";

	float var_1D_rrg(lat_times_lon);
	var_1D_rrg:long_name = "Variable for 2D irregular grid stored as 1D arrays";

	float var_2D_rct(lat,lon);
	var_2D_rct:long_name = "Variable for 2D rectangular grid stored as 2D array";

	float var_2D_rrg(lat,lon);
	var_2D_rrg:long_name = "Variable for 2D irregular grid stored as 2D array";

	float var_nm-dash;
	var_nm-dash:long_name = "Variable and attribute names include dash characters";
	var_nm-dash:att_nm-dash = 1.0e36f;

	float vld_rng(time);
	vld_rng:long_name = "Temperature";
	vld_rng:purpose = "Array containing _FillValue at some locations, out-of-range values at other locations, and valid data in the remainder";
	vld_rng:_FillValue = -999.0f;
	vld_rng:valid_min = 180.f;
	vld_rng:valid_max = 360.f;

//	float var_nm.dot;
//	var_nm.dot:long_name = "Variable and attribute names include dot characters";
//	20070102: Periods in attribute names choke OPeNDAP from FC7 RPM TODO nco911
//	20091105: Periods in attribute names choke ncgen   from RHEL5   TODO nco911
//	var_nm.dot:att_nm.dot = 1.0e36f;

	float wnd_spd(time,lat,lon);
	wnd_spd:long_name = "wind speed";
	wnd_spd:units = "meter second-1";
	wnd_spd:_FillValue = -999.0f;

data:
//	netCDF4-specific atomic types:
	int64_var_max=9223372036854775807;
	int64_var=73;
	string_var="If you prick us, do we not bleed? If you tickle us, do we not laugh? If you poison us, do we not die? And if you wrong us, shall we not revenge?";
	string_arr_var="20130723: Arrays of NC_STRING are simply separated by commas.","If there are commas within a string, well, then, be careful. Did we \"jump the shark\"?","This array comprises three sentences.","Woops, I mean four.";
         
	string_greek="alpha","beta","gamma","delta","epsilon","zeta","theta","iota"; 

	string_var2="20131121: This NC_STRING contains NCO's default XML string separator, *. And it contains multiple sequential copies of that separator, ***. Be sure ncks automatically switches to a different separator, aka the backup separator, the string obtained by removing the two spaces from this:\"* | *\". As of 20131121, ncks handles this correctly, yet toolsui breaks when trying to input the ncks-generated NcML. Appears to be a toolsui bug.";

	ubyte_var='z';
	uint_var_max=4294967295;
	uint_var=73;
//	uint64_var = 18446744073709551615; // 20131120: XML treats unsigned as signed types, so toolsui produces errors when reading maximum uint64 values (though not when reading maxium ubyte, ushort, and uint values)
	uint64_var=0;
	ushort_var=65535;

//	None in this file
//	netCDF3 atomic types:
	att_var=10.0,10.1,10.20,10.3000,10.40101,10.500001,10.60000001,10.7000001,10.80,10.9900;
	att_var_jsn=73;
	att_var_spc_chr=73;
	att_sng=20;
	area=10.,10.;
	area2=20.,5.;
	area_asm=1.,2.;
	areacella=1.,1.,2.,2.,3.,3.,4.,4.;
	bnd_var=1,2,3,4,5,6;
	byt_arr=0,1,2,3,4,5,6,7;
	byt_2D=0,1,2,3,4,5,6,7;
	byt_3D=0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23;
	byt_3D_rec= 	 1, 2, 3, 4, 5, 6, 7, 8,
			 9,10,11,12,13,14,15,16,
			17,18,19,20,21,22,23,24,
			25,26,27,28,29,30,31,32,
  			33,34,35,36,37,38,39,40,
			41,42,43,44,45,46,47,48,
			49,50,51,52,53,54,55,56,
			57,58,59,60,61,62,63,64,
			65,66,67,68,69,70,71,72,
			73,74,75,76,77,78,79,80;
	byt_bln_3D_rec=	0,0,0,0,0,0,0,0,
			0,0,0,0,0,0,0,1,
			0,0,0,0,0,0,1,1,
			0,0,0,0,0,1,1,1,
			0,0,0,0,1,1,1,1,
			0,0,0,1,1,1,1,1,
			0,0,1,1,1,1,1,1,
			0,1,1,1,1,1,1,1,
			1,1,1,1,1,1,1,1,
			1,0,1,0,1,0,1,0;

	byte_var='z';
	byte_var_neg=-122;
	char_var="z";
	// 20131015: This confuses the XML parser
	//	char_var_multinul="\b\n\0";
	// char_var_multinul='0','\n','\0';
	// 20180111: Historically we specified char_var_nul as '\0'
	// However, ncgen apparently turns '\0' into a zero
	// "correct" (meaning ncgen-supported) way to specify a scalar NUL character is with ""
	// As of today we specify char_var_nul as "" and char_var_nul_c_format as '\0'
	// char_var_nul_c_format indicates what happens when specifying characters in C-format
	// I think ncgen should support C-format byte codes for characters, though ncgen does not yet do so correctly
	char_var_nul="";
	char_var_nul_c_format='\0';
	char_var_zero="0";
	char_var_space=" ";
        char_var_1D_arr="two words";
        char_var_2D_arr="one","two";
        cnv_CF_grd=1,2,3,4,5,6,7,8;
	albers_conical_equal_area="";
	cnv_CF_crd=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8;
	cnv_CF_ncl=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	cnv_CF_ncl_var_1=11.,22.,23.,24.,25.,26.,27.,28.,29.,30.;
	cnv_CF_ncl_var_2=21.,32.,33.,34.,35.,36.,37.,38.,39.,40.;
	date_int=1964,3,12,12,9;
	dgn=73;
	dgn_var=73;
	double_var=10.;
	double_var2=10.;
	dps_dry=73;
	dps_wet=73;
	dps_ttl=73;
	e_dbl=2.71828182846;
	e_flt=2.71828182846;
// 	20100809: Single quotes around NC_CHAR coordinates required as of 4.1.2-beta1-snapshot2010080820
// 	20100809: Double quotes cause "String constant too long" error in ncgen
	fl_dmn='a','b','3';
	fl_nm="/home/zender/nco/data/in.cdl";
	float_var=10.;
	four=4.;
	g=9.8;
	grv_sfc=9.80665;
	vmr_CO2=400e-6;
	mmr_CO2=611e-6;
	gw=10.,10.;
	gw_T42=-87.863799,-85.096527,-82.312913,-79.525607,-76.736900,-73.947515,-71.157752,-68.367756,-65.577607,-62.787352,-59.997020,-57.206632,-54.416200,-51.625734,-48.835241,-46.044727,-43.254195,-40.463648,-37.673090,-34.882521,-32.091944,-29.301360,-26.510769,-23.720174,-20.929574,-18.138971,-15.348365,-12.557756,-9.767146,-6.976534,-4.185921,-1.395307,1.395307,4.185921,6.976534,9.767146,12.557756,15.348365,18.138971,20.929574,23.720174,26.510769,29.301360,32.091944,34.882521,37.673090,40.463648,43.254195,46.044727,48.835241,51.625734,54.416200,57.206632,59.997020,62.787352,65.577607,68.367756,71.157752,73.947515,76.736900,79.525607,82.312913,85.096527,87.863799;
	hyam=0.0036,0.0019894,0.0;
	hyai=0.002255,0.0438226,0.0,0.0;
	hybm=0.0,0.52,0.992;
	hybi=0.0,0.457453,0.985,1.0;
	P0=100000;
	gds_crd=0,1,2,3,4,5,6,7;
	gds_var=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8;
	gds_var_ncd=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8;
	gds_3dvar=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8,
	          274.1,274.2,274.3,274.4,274.5,274.6,274.7,274.8,
	          275.1,275.2,275.3,275.4,275.5,274.5,275.7,275.8,
	          276.1,276.2,276.3,276.4,276.5,276.5,276.7,276.8,
	          277.1,277.2,277.3,277.4,277.5,277.5,277.7,277.8,
	          278.1,278.2,278.3,278.4,278.5,278.6,278.7,278.8,
	          279.1,279.2,279.3,279.4,279.5,279.9,279.7,279.8,
	          280.1,280.2,280.3,280.4,280.5,280.9,280.7,280.8,
	          281.1,281.2,281.3,281.4,281.5,281.9,281.7,281.8,
	          282.1,282.2,282.3,282.4,282.5,282.9,282.7,282.8;
	lat_gds=-90, -30,  -30,    0,   0, 30,  30,  90;
	lon_gds=  0,   0,  180,    0, 180,  0, 180,   0;
	lat_gds_ncd=-90, -30,  -30,    0,   0, 30,  30,  90;
	lon_gds_ncd=  0,   0,  180,    0, 180,  0, 180,   0;
	lat=-90,90;
	lat_bnd=-90,0,0,90;
        lat_cal=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	lon_cal=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	lat_times_lon=0,1,2,3,4,5,6,7;
	lat_times_lon_nbr=8;
	lat_1D_rct=-90, -90,  -90,  -90,  90, 90,  90,  90;
	lon_1D_rct=  0,  90,  180,  270,   0, 90, 180, 270;
	lat_1D_rrg=-90, -30,  -30,    0,   0, 30,  30,  90;
	lon_1D_rrg=  0,   0,  180,    0, 180,  0, 180,   0;
	lat_2D_rct=-90, -90,  -90,  -90,  90, 90,  90,  90;
	lon_2D_rct=  0,  90,  180,  270,   0, 90, 180, 270;
	lat_2D_rrg=-90, -30,  -30,    0,   0, 30,  30,  90;
	lon_2D_rrg=  0,   0,  180,    0, 180,  0, 180,   0;
	lat_grd=-90,0,90;
	lat_cpy=-90,90;
	lat_var=1.,2.;
	lat_wgt=1.,2.;
//	lat_T42=0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63;
	lat_T42=-88.240089,-85.092445,-82.311981,-79.525253,-76.736732,-73.947418,-71.157700,-68.367722,-65.577576,-62.787331,-59.997005,-57.206619,-54.416191,-51.625729,-48.835236,-46.044724,-43.254192,-40.463646,-37.673088,-34.882519,-32.091942,-29.301357,-26.510769,-23.720173,-20.929573,-18.138969,-15.348364,-12.557755,-9.767145,-6.976533,-4.185921,-1.395307,1.395307,4.185921,6.976533,9.767145,12.557755,15.348364,18.138969,20.929573,23.720173,26.510769,29.301357,32.091942,34.882519,37.673088,40.463646,43.254192,46.044724,48.835236,51.625729,54.416191,57.206619,59.997005,62.787331,65.577576,68.367722,71.157700,73.947418,76.736732,79.525253,82.311981,85.092445,88.240089;
	lsmlev=0.05,0.1,0.2,0.5,1.0,3.0;
	lev=100,500,1000;
	ilev=50,200,750,1005;
	lev_bnd=0,300,300,750,750,1013.25;
	lev_cpy=100,500,1000;
	lev_var=100.,500.,1000.;
	lev_wgt=10,2,1;
	lon=0,90,180,270;
	Lon=-180,-90,0,90;
	Lat=-45,45;
	LatLon=0,1,2,3,4,5,6,7;
	lond=0,90,180,270;
	lonf=0,90,180,270;
	lon_grd=-45,45,135,225,315;
	lon_wgt=0.347855,0.652145,0.652145,0.347855;
//	lon_T42=0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127;
	lon_T42=0.000000,2.812500,5.625000,8.437500,11.250000,14.062500,16.875000,19.687500,22.500000,25.312500,28.125000,30.937500,33.750000,36.562500,39.375000,42.187500,45.000000,47.812500,50.625000,53.437500,56.250000,59.062500,61.875000,64.687500,67.500000,70.312500,73.125000,75.937500,78.750000,81.562500,84.375000,87.187500,90.000000,92.812500,95.625000,98.437500,101.250000,104.062500,106.875000,109.687500,112.500000,115.312500,118.125000,120.937500,123.750000,126.562500,129.375000,132.187500,135.000000,137.812500,140.625000,143.437500,146.250000,149.062500,151.875000,154.687500,157.500000,160.312500,163.125000,165.937500,168.750000,171.562500,174.375000,177.187500,180.000000,182.812500,185.625000,188.437500,191.250000,194.062500,196.875000,199.687500,202.500000,205.312500,208.125000,210.937500,213.750000,216.562500,219.375000,222.187500,225.000000,227.812500,230.625000,233.437500,236.250000,239.062500,241.875000,244.687500,247.500000,250.312500,253.125000,255.937500,258.750000,261.562500,264.375000,267.187500,270.000000,272.812500,275.625000,278.437500,281.250000,284.062500,286.875000,289.687500,292.500000,295.312500,298.125000,300.937500,303.750000,306.562500,309.375000,312.187500,315.000000,317.812500,320.625000,323.437500,326.250000,329.062500,331.875000,334.687500,337.500000,340.312500,343.125000,345.937500,348.750000,351.562500,354.375000,357.187500;
	ppc_flt_2D=    -1,-2,-3,-4,-5,-6,-7,-8,-9,-10,
	               -11,-12,-13,-14,-15,-16,-17,-18,-19,-20;
	ppc_dbl=0.0,0.1,0.12,0.123,0.1234,0.12345,0.123456,0.1234567,0.12345678,0.123456789;
	ppc_flt=0.0,0.1,0.12,0.123,0.1234,0.12345,0.123456,0.1234567,0.12345678,0.123456789;
	ppc_big=123456789e-10,123456789e-9,123456789e-8,123456789e-7,123456789e-6,123456789e-5,123456789e-4,123456789e-3,123456789e-2,123456789e-1;
	ppc_btg=1234567890e20,1234567890e19,1234567890e18,1234567890e17,1234567890e16,1234567890e15,1234567890e14,1234567890e13,1234567890e12,1234567890e11;
	ppc_btg_scl=1234567890e11;
	ppc_hgh=0.00000000000000000000,0.10000000000000000000,0.12000000000000000000,0.123000000000000000000,0.1234000000000000000,0.12345000000000000000,0.123456000000000000000000,0.12345670000000000000000000,0.123456780000000000000,0.123456789000000000000;
	// 20220731 NCZarr I/O chokes here, apparently ncgen parses 15+ digit mantissas as integers? 20220819 that problem was fixed sometime before today, extended decimals now work fine
	ppc_hgr=0.123456789000000000000,0.1234567890100000000000,0.1234567890120000000000,0.12345678901230000000000,0.123456789012340000000,0.12345678901234500000,0.12345678901234560000,0.12345678901234567000,0.12345678901234567800,0.12345678901234567890;
        ppc_dcm=55,155,255,355,455,555,655,755,855,955;
        ppc_tst=0.0,_,0.1234567,-0.1234567,64,-64,123456789e25,123456789e-25,3.1415926535897932384626433832795029,-3.1415926535897932384626433832795029;
	ppc_zro_flt=0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0;
	ppc_zro_dbl=0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0;
	ppc_zro_int=0,0,0,0,0,0,0,0,0,0;
	qnt_flt_tst1=1.1111111;
	qnt_dbl_tst1=1.111111111111;
	qnt_flt_tst2=1.11111111, 1.0, 9.99999999, 12345.67, .1234567;
	// 20220731 NCZarr I/O chokes here, apparently ncgen parses 15+ digit mantissas as integers? 20220819 that problem was fixed sometime before today, extended decimals now work fine
	qnt_dbl_tst2=1.1111111, 1.0, 9.999999999, 1234567890.12345, 123456789012345.0;
	var_msk=0.,1.,0.,0.,1.,1.,0.,2.;
	var_mss_nil=0.,1.,2.,3.;
	var_mss_0=_,1.,2.,3.;
	var_mss_1=0.,_,2.,3.;
	var_mss_2=0.,1.,_,3.;
	var_mss_3=0.,1.,2.,_;
	ORO=0.,1.,0.,0.,1.,1.,0.,2.;
	orog=0.,1.,0.,0.,1.,1.,0.,2.;
	orog2=1.,1.,1.,1.,1.,1.,1.,1.;
	orog3=0.,0.,0.,0.,1.,1.,1.,1.;
	mask=0.,1.,0.,0.,1.,1.,0.,1.;
//	mask=0.,0.,0.,0.,0.,0.,0.,0.;
//	mask=1.,1.,1.,1.,1.,1.,1.,1.;
	fll_val=73,-999,73,-999;
	fll_val_mss_val=73,-999,73,-999;
	md5_a="a";
	md5_abc="abc";
	msk_prt_mss_prt=0.5,1.0e36,1.5,1.0e36;
	mss_val=73,1.0e36,73,1.0e36;
	mss_val_all=1.0e36,1.0e36,1.0e36,1.0e36;
	mss_val_fst=-999,73,-999,73;
	mss_val_scl=1.0e36;
	mss_val_scl_sml=1.0e4;
	//nan_arr=0,nan;
	nan_arr=0,73;
	//nan_scl=nan;
	nan_scl=1;
	negative_one=-1.;
	nm_pnd=1;
	nm_spc=1;
	no_mss_val=73,1.0e36,73,1.0e36;
	non_nul_trm_char_one_dmn='a','b';
	non_nul_trm_char_two_dmn="abcd","efgh","ijkm";
	one=1.;
	one_dmn_rec_var=1,2,3,4,5,6,7,8,9,10;
	one_dmn_rec_wgt=2,1,0,0,0,0,0,0,0,0;
	one_dmn_rec_var_unsorted=10,4,6,2,8,1,9,7,3,5;
	one_dmn_rec_var_flt=1,2,3,4,5,6,7,8,9,10;
	one_dmn_rec_var_flt_mss=_,2,3,4,5,6,7,8,9,_;
	one_dmn_rec_var_flt_scl=1,2,3,4,5,6,7,8,9,10;
// First use of underscore to indicate _FillValue in in.cdl is here in one_dmn_rec_var_flt_mss_scl on 20140916
	one_dmn_rec_var_flt_mss_scl=_,2,3,4,5,6,7,8,9,_;
	one_dmn_rec_var_dbl=1,2,3,4,5,6,7,8,9,10;
	one_dmn_rec_var_missing_value=1,2,3,4,5,6,7,8,9,1.0e36;
	one_dmn_rec_var_mss_val=1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36;
	one_dmn_rec_var_mss_val_arr=1,2,3,4,5,6,7,8,9,10;
	one_dmn_rec_var__FillValue=1,2,3,4,5,6,7,8,9,1.0e36;
	one_dmn_rec_var_unsorted__FillValue=1.0e36,4,6,2,8,1,9,7,3,5;
	one_dmn_rec_var_mdn=1,1,2,2,2,2,10,10,10,10;
	one_dmn_rec_var_mdn__FillValue=1,-999,2,2,-999,-999,10,10,10,-999;
	RDM=1,9,36,84,126,126,84,36,9,1;
	one_dmn_rec_var_sng="Hello Worl";
	one_dmn_var=1.,10.;
	one_dmn_int_val_one=1,1;
	one_dmn_int_val_two=2,2;
	pck=1;
	pck_3=1;
	pck_5=2;
	pck_7=1;
	rec_var_pck_scale_factor_only=1,2,3,4,5,6,7,8,9,10;
	pck_arr=-32767,0,1,32767;
	pck_crd=-32767,0,1,32767;
	pi=3.1415926535897932384626433832795029;
	pi1=3.1415927,3.1415937,3.1415946,3.1415956,3.1415966,3.1415977,3.1415987,3.1415997,3.1416006,3.1416016;
	pi2=3.1415927,3.1415937,3.1415946,3.1415956,3.1415966,3.1415977,3.1415987,3.1415997,3.1416006,3.1416016;
	pi3=3.1415927,3.1415937,3.1415946,3.1415956,3.1415966,3.1415977,3.1415987,3.1415997,3.1416006,3.1416016;
	pi4=3.1415927,3.1415937,3.1415946,3.1415956,3.1415966,3.1415977,3.1415987,3.1415997,3.1416006,3.1416016;
	pi5=3.1415927,3.1415937,3.1415946,3.1415956,3.1415966,3.1415977,3.1415987,3.1415997,3.1416006,3.1416016;
	pi6=3.1415927,3.1415937,3.1415946,3.1415956,3.1415966,3.1415977,3.1415987,3.1415997,3.1416006,3.1416016;
	pi7=3.1415927,3.1415937,3.1415946,3.1415956,3.1415966,3.1415977,3.1415987,3.1415997,3.1416006,3.1416016;
	pi_arr_dbl=3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029;
	pi_arr_flt=3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029,3.1415926535897932384626433832795029;
	upk=3.;
	upk_arr=-32767.,0.,1.,32767.;
	H2O=1.0;
	H2OH2O=1.0;
	H2SO4=1.0;
	H2O_lqd=1.0;
	H2O_ice=1.0;
	Q=1.0e36;
	Q1=1.0e36;
	AQ01=1.0e36;
	QQ01=1.0e36;
	QA01=1.0e36;
	Q01Q=1.0e36;
	Q01=1;
	Q02=2;
	Q03=3;
	Q04=4;
	Q05=5;
	Q06=6;
	Q07=7;
	Q08=8;
	Q09=9;
	Q10=10;
	Q11=11;
	Q12=12;
	Q13=13;
	Q14=14;
	Q15=15;
	Q16=16;
	Q17=17;
	Q18=18;
	Q19=19;
	Q20=20;
	Q21=21;
	Q22=22;
	Q23=23;
	Q24=24;
	Q25=25;
	Q26=26;
	Q27=27;
	Q28=28;
	Q29=29;
	Q30=30;
	Q31=31;
	Q32=32;
	Q33=33;
	Q34=34;
	Q35=35;
	Q36=36;
	Q37=37;
	Q38=38;
	Q39=39;
	Q40=40;
	Q41=41;
	Q42=42;
	Q43=43;
	Q44=44;
	Q45=45;
	Q46=46;
	Q47=47;
	Q48=48;
	Q49=49;
	Q50=50;
	Q51=51;
	Q52=52;
	Q53=53;
	Q54=54;
	Q55=55;
	Q56=56;
	Q57=57;
	Q58=58;
	Q59=59;
	Q60=60;
	Q61=61;
	Q62=62;
	Q63=63;
	Q64=64;
	Q65=65;
	Q66=66;
	Q67=67;
	Q68=68;
	Q69=69;
	Q70=70;
	Q71=71;
	Q72=72;
	Q73=73;
	Q74=74;
	Q75=75;
	Q76=76;
	Q77=77;
	Q78=78;
	Q79=79;
	Q80=80;
	Q81=81;
	Q82=82;
	Q83=83;
	Q84=84;
	Q85=85;
	Q86=86;
	Q87=87;
	Q88=88;
	Q89=89;
	Q90=90;
	Q91=91;
	Q92=92;
	Q93=93;
	Q94=94;
	Q95=95;
	Q96=96;
	Q97=97;
	Q98=98;
	Q99=99;
	Q100=100;
	non_rec_var_flt_pck=1,2,3,4;
	rec_var_dbl=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	rec_var_dbl_mss_val_dbl_pck=-999,32767,21845,10922,0,-10922,-21845,-32767,-999,-999;
	rec_var_dbl_mss_val_dbl_pck_lng=-999,32767,21845,10922,0,-10922,-21845,-32767,-999,-999;
	rec_var_dbl_mss_val_sht_pck_sht=-999,32767,21845,10922,0,-10922,-21845,-32767,-999,-999;
	rec_var_flt_mss_val_flt_pck_flt=-9.96921e+33,0.032,0.033,0.034,0.035,0.036,0.037,0.038,-9.96921e+33,-9.96921e+33;
	SALT=-9.96921e+33,0.032,0.033,0.034,0.035,0.036,0.037,0.038,-9.96921e+33,-9.96921e+33;
	rec_var_dbl_mss_val_dbl_upk=-999.,2.,3.,4.,5.,6.,7.,8.,-999.,-999.;
	rec_var_dbl_mss_val_sht_pck=-999,32767,21845,10922,0,-10922,-21845,-32767,-999,-999;
	rec_var_dbl_mss_val_sht_upk=-999.,2.,3.,4.,5.,6.,7.,8.,-999.,-999.;
	rec_var_dbl_pck=1,2,3,4,5,6,7,8,9,10;
	rec_var_flt=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	rec_var_flt_mss_val_dbl=1.0e36,2.,3.,4.,5.,6.,7.,8.,1.0e36,1.0e36;
	rec_var_flt_mss_val_flt=1.0e36,2.,3.,4.,5.,6.,7.,8.,1.0e36,1.0e36;
	rec_var_flt_mss_val_flt_all=1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36;
	rec_var_flt_mss_val_flt_all_but_one=1.0e36,1.0e36,1.0e36,1.0e36,5.0,1.0e36,1.0e36,1.0e36,1.0e36,1.0e36;
	rec_var_flt_mss_val_flt_all_but_two=1.0e36,1.0e36,1.0e36,1.0e36,5.0,1.0e36,1.0e36,1.0e36,1.0e36,10.0;
	rec_var_flt_mss_val_int=-999.,2.,3.,4.,5.,6.,7.,8.,-999.,-999.;
	rec_var_flt_pck=1,2,3,4,5,6,7,8,9,10;
	rec_var_int_mss_val_dbl=-999,2,3,4,5,6,7,8,-999,-999;
	rec_var_int_mss_val_flt=-999,2,3,4,5,6,7,8,-999,-999;
	rec_var_int_mss_val_int=-999,2,3,4,5,6,7,8,-999,-999;
	rlev=1000,500,100;
	rz=0,5000,17000;
	scl_dbl_pck=10922;
	scalar_var=10.;
	short_var=10;
	three=3.;
	three_dmn_var=0.,1.,2.,3.,4.,5.,6.,7.,8.,9.,10.,11.,12.,13.,14.,15.,16.,17.,18.,19.,20.,21.,22.,23.;
	three_dmn_var_crd=0.,1.,2.,3.,12.,13.,14.,15.,4.,5.,6.,7.,16.,17.,18.,19.,8.,9.,10.,11.,20.,21.,22.,23.;
	three_dmn_var_cf=0.,1.,2.,3.,12.,13.,14.,15.,4.,5.,6.,7.,16.,17.,18.,19.,8.,9.,10.,11.,20.,21.,22.,23.;
	three_dmn_var_cf2=0.,1.,2.,3.,12.,13.,14.,15.,4.,5.,6.,7.,16.,17.,18.,19.,8.,9.,10.,11.,20.,21.,22.,23.;
	time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
        time_rpt=1.,2.,3.,1.,2.,3.,1.,2.,3.,1.;
	time_bnds=0.5,1.5,1.5,2.5,2.5,3.5,3.5,4.5,4.5,5.5,5.5,6.5,6.5,7.5,7.5,8.5,8.5,9.5,9.5,10.5;
	climatology_bounds=0.5,1.5,1.5,2.5,2.5,3.5,3.5,4.5,4.5,5.5,5.5,6.5,6.5,7.5,7.5,8.5,8.5,9.5,9.5,10.5;
	tm_scn=59;
	tm_std=59;
	tm_grg=59;
	tm_jln=59;
	tm_360=59;
	tm_365=59;
	tm_366=59;
	od=20,22,24,26,28,30,32,34,36,38;
	tpt=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8,273.9,274.0;
	tpt_flt=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8,273.9,274.0;
	tpt_dbl=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8,273.9,274.0;
	two=2.;
	two_dmn_var=1.5,5.5,9.5,13.5,17.5,21.5;
	u=1.,0.,1.,0.,1.,0.,1.,0.,1.,0.;
	v=0.,1.,0.,1.,0.,1.,0.,1.,0.,1.;
	val_half=0.5;
	val_half_half=0.5,0.5;
	val_max_max_sht=17000,17000;
	val_eminusten=1.1e-10;
	val_one_int=1;
	val_one_mss=1.,1.0e36;
	val_one_mss_int=1,-99;
	val_one_one_int=1,1;
	var_nm-dash=1.0;
//	var_nm.dot=1.0;
	var_1D_rct=0.,1.,0.,0.,1.,1.,0.,2.;
	var_1D_rrg=0.,1.,0.,0.,1.,1.,0.,2.;
	var_2D_rct=0.,1.,0.,0.,1.,1.,0.,2.;
	var_2D_rrg=0.,1.,0.,0.,1.,1.,0.,2.;
	weight=10.,10.;
	wgt_one=1.,1.;
	wvl=0.5e-6,1.0e-6;
	z=17000,5000,0;
	zero=0.;
// 	        date=640312,640313,640314,640315,640316,640317,640318,640319,640320,640321;
	date=640224,640225,640226,640227,640228,640301,640302,640303,640304,640305;
 	int_var=10;
 	long_var=10;
 	nbdate=640224;
	fl_nm_arr="/data/zender/dstccm04/dstccm04_8589_01.nc",
		"/data/zender/dstccm04/dstccm04_8589_02.nc",
		"/data/zender/dstccm04/dstccm04_8589_03.nc";
	fl_nm_rec="/data/zender/dstccm04/dstccm04_8589_01.nc",
	  "/data/zender/dstccm04/dstccm04_8589_02.nc",
	  "/data/zender/dstccm04/dstccm04_8589_03.nc",
	  "/data/zender/dstccm04/dstccm04_8589_04.nc",
	  "/data/zender/dstccm04/dstccm04_8589_05.nc",
	  "/data/zender/dstccm04/dstccm04_8589_06.nc",
	  "/data/zender/dstccm04/dstccm04_8589_07.nc",
	  "/data/zender/dstccm04/dstccm04_8589_08.nc",
	  "/data/zender/dstccm04/dstccm04_8589_09.nc",
	  "/data/zender/dstccm04/dstccm04_8589_10.nc";
	date_sng="2010-11-01T00:00:00.000000";
	date_rec="2010-11-01T00:00:00.000000",
	  "2010-11-01T01:00:00.000000",
	  "2010-11-01T02:00:00.000000",
	  "2010-11-01T03:00:00.000000",
	  "2010-11-01T04:00:00.000000",
	  "2010-11-01T05:00:00.000000",
	  "2010-11-01T06:00:00.000000",
	  "2010-11-01T07:00:00.000000",
	  "2010-11-01T08:00:00.000000",
	  "2010-11-01T09:00:00.000000";
	time_lon=0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0;
	two_dmn_rec_var_sng="abc",
				"bcd",
				"cde",
				"def",
				"efg",
				"fgh",
				"ghi",
				"hij",
				"jkl",
				"klm";
	two_dmn_rec_var=1.,2.0,3.,
			1.,2.1,3.,
			1.,2.2,3.,
			1.,2.3,3.,
			1.,2.4,3.,
			1.,2.5,3.,
			1.,2.6,3.,
			1.,2.7,3.,
			1.,2.8,3.,
			1.,2.9,3.;
	three_dmn_rec_var= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
  				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				73,74,75,76,77,78,79,80;
	three_dmn_rec_var_pck=  32766, 31936, 31107, 30277, 29448, 28618, 27789, 26959, 
	  26130, 25300, 24471, 23641, 22812, 21982, 21153, 20323, 
	  19494, 18664, 17835, 17005, 16176, 15346, 14517, 13687, 
	  12858, 12028, 11199, 10369, 9539, 8710, 7880, 7051, 
	  6221, 5392, 4562, 3733, 2903, 2074, 1244, 415, 
	  -415, -1244, -2074, -2903, -3733, -4562, -5392, -6221, 
	  -7051, -7880, -8710, -9539, -10369, -11199, -12028, -12858, 
	  -13687, -14517, -15346, -16176, -17005, -17835, -18664, -19494, 
	  -20323, -21153, -21982, -22812, -23641, -24471, -25300, -26130, 
	  -26959, -27789, -28618, -29448, -30277, -31107, -31936, -32766 ; 
	prs_sfc=		 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
  				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				73,74,75,76,77,78,79,80;
	PS=			101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
  				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325,
				101325,101325,101325,101325,101325,101325,101325,101325;
	three_dmn_var_dbl= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				-99,-99,-99,-99,-99,-99,-99,-99,
				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				-99,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				-99,74,75,76,77,78,79,-99;
	zg=              	 1, 2, 3, 4, 5, 6, 7, 8,9,10,11,12,
				13,14,15,16,17,18,19,20,21,22,23,24,
	                        25,26,27,28,29,30,31,32,33,34,35,36,
				37,38,39,40,41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,57,58,59,60,
                                61,62,63,64,65,66,67,68,69,70,71,72,
				73,74,75,76,77,78,79,80,81,82,83,84,
                                85,86,87,88,89,90,91,92,93,94,95,96,
                                97,98,99,100,101,102,103,104,105,106,107,108,
                                109,110,111,112,113,114,115,116,117,118,119,120;
	three_dmn_var_int= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				-99,-99,-99,-99,-99,-99,-99,-99,
				25,26,27,28,29,30,31,32,
				33,34,35,36,37,38,39,40,
				41,-99,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				-99,58,59,60,-99,62,63,64,
				65,-99,67,68,69,70,71,72,
				-99,74,75,-99,77,78,79,80;
	three_dmn_var_sht= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 -99,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
				-99,34,35,-99,37,38,39,40,
				41,42,43,44,-99,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,-99,61,62,63,64,
				65,66,67,68,69,70,71,72,
				-99,-99,-99,-99,-99,-99,-99,-99;
	th=			1, 2, 3, 4, 5, 6, 7, 8,
				9,10,11,12,13,14,15,16,
			  	17,18,19,20,21,22,23,24,
			  	-99,-99,-99,-99,-99,-99,-99,-99,
			  	33,34,35,36,37,38,39,40,
			  	41,42,43,44,45,46,47,48,
			  	49,50,51,52,53,54,55,56,
			  	-99,58,59,60,61,62,63,64,
			  	65,66,67,68,69,70,71,72,
			 	-99,74,75,76,77,78,79,-99;
	four_dmn_rec_var= 	  1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12,
				 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24,
				 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36,
				 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48,
				 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60,
				 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72,
				 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84,
				 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96,
				 97, 98, 99,100,101,102,103,104,105,106,107,108,
				109,110,111,112,113,114,115,116,117,118,119,120,
				121,122,123,124,125,126,127,128,129,130,131,132,
				133,134,135,136,137,138,139,140,141,142,143,144,
				145,146,147,148,149,150,151,152,153,154,155,156,
				157,158,159,160,161,162,163,164,165,166,167,168,
				169,170,171,172,173,174,175,176,177,178,179,180,
				181,182,183,184,185,186,187,188,189,190,191,192,
				193,194,195,196,197,198,199,200,201,202,203,204,
				205,206,207,208,209,210,211,212,213,214,215,216,
				217,218,219,220,221,222,223,224,225,226,227,228,
				229,230,231,232,233,234,235,236,237,238,239,240;
	td=		1,2,3,4,5,6,7,8,9,10;
	tx=		1,2,3,4,5,6,7,8,9,10,
			11,12,13,14,15,16,17,18,19,20,
			21,22,23,24,25,26,27,28,29,30,
			31,32,33,34,35,36,37,38,39,40;
	ty=		1,2,3,4,5,6,7,8,9,10,
			11,12,13,14,15,16,17,18,19,20;
	tz=		1,2,3,4,5,6,7,8,9,10,
			11,12,13,14,15,16,17,18,19,20,
			21,22,23,24,25,26,27,28,29,30;
	tyz=		1,2,3,4,5,6,7,8,9,10,
			11,12,13,14,15,16,17,18,19,20,
			21,22,23,24,25,26,27,28,29,30,
	                31,32,33,34,35,36,37,38,39,40,
                        41,42,43,44,45,46,47,48,49,50,
			51,52,53,54,55,56,57,58,59,60;
	xyz=0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23;
	txyz=		 	  1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12,
				 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24,
				 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36,
				 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48,
				 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60,
				 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72,
				 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84,
				 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96,
				 97, 98, 99,100,101,102,103,104,105,106,107,108,
				109,110,111,112,113,114,115,116,117,118,119,120,
				121,122,123,124,125,126,127,128,129,130,131,132,
				133,134,135,136,137,138,139,140,141,142,143,144,
				145,146,147,148,149,150,151,152,153,154,155,156,
				157,158,159,160,161,162,163,164,165,166,167,168,
				169,170,171,172,173,174,175,176,177,178,179,180,
				181,182,183,184,185,186,187,188,189,190,191,192,
				193,194,195,196,197,198,199,200,201,202,203,204,
				205,206,207,208,209,210,211,212,213,214,215,216,
				217,218,219,220,221,222,223,224,225,226,227,228,
				229,230,231,232,233,234,235,236,237,238,239,240;

//	three_double_dmn= 	 1, 2, 3, 4, 5, 6, 7, 8,
//				 9,10,11,12,13,14,15,16,
//				17,18,19,20,21,22,23,24,
//				-99,-99,-99,-99,-99,-99,-99,-99,
//				33,34,35,36,37,38,39,40,
//				41,42,43,44,45,46,47,48,
//				49,50,51,52,53,54,55,56,
//				-99,58,59,60,61,62,63,64,
//				65,66,67,68,69,70,71,72,
//				-99,74,75,76,77,78,79,-99,
//				1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5,
//				 9.5,10.5,11.5,12.5,13.5,14.5,15.5,16.5,
//				17.5,18.5,19.5,20.5,21.5,22.5,23.5,24.5,
//				-99.5,-99.5,-99.5,-99.5,-99.5,-99.5,-99.5,-99.5,
//				33.5,34.5,35.5,36.5,37.5,38.5,39.5,40.5,
//				41.5,42.5,43.5,44.5,45.5,46.5,47.5,48.5,
//				49.5,50.5,51.5,52.5,53.5,54.5,55.5,56.5,
//				-99.5,58.5,59.5,60.5,61.5,62.5,63.5,64.5,
//				65.5,66.5,67.5,68.5,69.5,70.5,71.5,72.5,
//				-99.5,74.5,75.5,76.5,77.5,78.5,79.5,-99.5;
				
        time_int_udunits = 86400;

	time_udunits = 876012, 876018, 876024;

	vld_rng=		273.,-999.,180.,179.,273.,360.,361.,1.0e36,-1.0e36,273.;

	wnd_spd=		-999,0.5,1.5,0.5,1.5,0.5,1.5,0.5,
				0.5,-999,0.5,0.5,0.5,0.5,0.5,0.5,
				0.5,1.5,-999,1.5,0.5,1.5,0.5,1.5,
				0.5,0.5,0.5,-999,0.5,0.5,0.5,0.5,
  				1.5,1.5,1.5,1.5,-999,1.5,1.5,1.5,
				0.5,0.5,0.5,0.5,0.5,-999,0.5,0.5,
				2.5,2.5,2.5,2.5,2.5,2.5,-999,2.5,
				0.5,0.5,0.5,0.5,0.5,0.5,0.5,-999,
				0.5,0.5,0.5,0.5,0.5,0.5,0.5,0.5,
				0.5,0.5,2.5,0.5,0.5,2.5,0.5,0.5;
} // end netcdf







