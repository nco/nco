// Generate netCDF file with:
// ncgen -k netCDF-4 -b -o ~/nco/data/cmip5.nc ~/nco/data/cmip5.cdl

netcdf cmip5 {
  dimensions:
  time=unlimited;
 
  //
  //cesm
  //
  group: cesm { 
  variables:
  float tas(time);
  data:
  tas=272,272,272,272;
  } // end cesm
  
  //
  //ecmwf
  //
  group: ecmwf { 
  variables:
  float tas(time);
  data:
  tas=273,273,273,273;
  } // end ecmwf
  
  //
  //gfdl
  //
  group: gfdl { 
  variables:
  float tas(time);
  data:
  tas=274,274,274,274;
  } // end gfdl

} // end root group
