// Purpose: CDL file to generate netCDF test file

// Usage:
// ncgen -b -o in.nc in.cdl
// ncgen -b -o /home/zender/nc/nco/data/in.nc /home/zender/nc/nco/data/in.cdl
// mswrite -t 365 in.nc /ZENDER/tmp/in.nc
// mswrite -t 365 in.nc /ZENDER/tmp/h0001.nc
// mswrite -t 365 in.nc /ZENDER/tmp/h0002.nc
// mswrite -t 365 in.nc /ZENDER/tmp/h0003.nc
// mswrite -t 365 in.nc /ZENDER/tmp/h0004.nc

// NB: Changing the values of the variables below, especially the coordinate 
// variables, may affect the outcome of the test script nco_tst.sh.

// NCL usage:
// id_in=addfile("/home/zender/nc/nco/data/in.nc","r")
// print(id_in)
// list_filevars(id_in)

netcdf in {
dimensions:
	band=2,lat=2,lev=3,rlev=3,lon=4,time=unlimited;
variables:
	:convention = "NCAR-CSM";
	:history = "History global attribute.\n";
	:julian_day = 200000.04;
	:RCS_Header = "$Header: /data/zender/nco_20150216/nco/data/in.cdl,v 1.7 1999-05-11 08:01:06 zender Exp $";

	float lat(lat);
	float lat_var(lat);
	float lat_wgt(lat);
	float lev(lev);
	lev:purpose = "Monotonically increasing coordinate pressure";
	float rlev(rlev);
	rlev:purpose = "Monotonically decreasing coordinate pressure";
	float lon(lon);
	double time(time);

	long nbdate;
	nbdate:long_name = "base date as 6 or 8 digit integer (YYMMDD or YYYYMMDD)";
	long date(time);
	date:long_name = "current date as 6 or 8 digit integer (YYMMDD or YYYYMMDD)";

	float mss_val(lon);
	mss_val:long_name = "missing value example";
	mss_val:missing_value = 1.0e36f;

	float no_mss_val(lon);
	no_mss_val:long_name = "no missing value";

	float scalar_var;
	scalar_var:long_name = "scalar variable";
	scalar_var:units = "Fraction";

	float float_var;
	float_var:long_name = "float";

	double double_var;
	double_var:long_name = "double";

	long long_var;
	long_var:long_name = "long";

	short short_var;
	short_var:long_name = "short";

	char char_var;
	char_var:long_name = "char";

	byte byte_var;
	byte_var:long_name = "byte";

	float zero;
	zero:long_name = "zero";

	float one;
	one:long_name = "one";

	float two;
	two:long_name = "two";

	float three;
	three:long_name = "three";

	float negative_one;
	negative_one:long_name = "negative one";

	float lev_var(lev);
	lev_var:long_name = "lev_var";

	float lev_wgt(lev);
	lev_wgt:long_name = "lev_wgt";

	float g;
	g:long_name = "g";

	float z(lev);
	z:long_name = "Height";
	z:units = "meter";
	z:purpose = "Height stored with a monotonically increasing coordinate";

	float rz(rlev);
	rz:long_name = "Height";
	rz:units = "meter";
	rz:purpose = "Height stored with a monotonically decreasing coordinate";

	float one_dim_var(band);

	float att_var;
	att_var:byte_att = '\0';
	att_var:char_att = "Sentence one.\nSentence two.\n";
	att_var:short_att = 37s;
	att_var:long_att = 73l;
	att_var:float_att = 73.f,72.f,71.f;
	att_var:double_att = 73.d;

	long band_var(lev,band);
	band_var:byte_att = '\0';
	band_var:char_att = "Sentence one.\nSentence two.\n";
	band_var:short_att = 37s;
	band_var:long_att = 73l;
	band_var:float_att = 73.f;
	band_var:double_att = 73.d;

	float three_dim_var(lat,lev,lon);
	three_dim_var:long_name = "three dimensional variable";
	three_dim_var:units = "Fraction";

	float two_dim_var(lat,lev);
	two_dim_var:long_name = "two dimensional variable";
	two_dim_var:units = "Fraction";

	float mask(lat,lon);
	mask:long_name = "mask variable like ORO";
	mask:units = "Fraction";

	float ORO(lat,lon);
	ORO:long_name = "Orography";
	ORO:units = "Fraction";

	float weight(lat);
	weight:long_name = "Gaussian weight";
	weight:units = "Fraction";

	float gw(lat);
	gw:long_name = "gw variable like gw";
	gw:units = "Fraction";

	float rec_var_flt(time);
	rec_var_flt:long_name = "record variable, float";

	double rec_var_dbl(time);
	rec_var_dbl:long_name = "record variable, double";

	long one_dim_rec_var(time);
	one_dim_rec_var:long_name = "one dimensional record variable";
	one_dim_rec_var:units = "second";

	char one_dim_rec_var_sng(time);
	one_dim_rec_var_sng:long_name = "one dimensional record variable of string";

	char two_dim_rec_var_sng(time,lev);
	two_dim_rec_var_sng:long_name = "two dimensional record variable of string";

	float two_dim_rec_var(time,lev);
	two_dim_rec_var:long_name = "two dimensional record variable";
	two_dim_rec_var:units = "watt meter-2";

	float three_dim_rec_var(time,lat,lon);
	three_dim_rec_var:long_name = "three dimensional record variable";
	three_dim_rec_var:units = "watt meter-2";

	float four_dim_rec_var(time,lat,lev,lon);
	four_dim_rec_var:long_name = "four dimensional record variable";
	four_dim_rec_var:units = "watt meter-2";

data:
	lat=-90,90;
	lev=100,500,1000;
	rlev=1000,500,100;
	lon=0,90,180,270;
	time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	mss_val=73,1.0e36,73,1.0e36;
	no_mss_val=73,1.0e36,73,1.0e36;
	scalar_var=10.;
	att_var=10.;
	lat_var=1.,2.;
	lat_wgt=1.,2.;
	lev_var=100.,500.,1000.;
	lev_wgt=10,2,1;
	zero=0.;
	one=1.;
	two=2.;
	three=3.;
	negative_one=-1.;
	g=9.8;
 	nbdate=640312;
 	date=640312,640313,640314,640315,640316,640317,640318,640319,640320,640321;
	float_var=10.;
	double_var=10.;
	short_var=10;
 	long_var=10;
	char_var="z";
	byte_var='z';
	one_dim_var=1.,10.;
	z=17000,5000,0;
	rz=0,5000,17000;
	band_var=1,2,3,4,5,6;
	two_dim_var=1.5,5.5,9.5,13.5,17.5,21.5;
	weight=10.,10.;
	gw=10.,10.;
	ORO=1.,1.,1.,1.,1.,1.,1.,1.;
	mask=0.,1.,0.,0.,1.,1.,0.,2.;
//	mask=1.,1.,1.,1.,1.,1.,1.,1.;
//	mask=0.,0.,0.,0.,0.,0.,0.,0.;
	three_dim_var=0.,1.,2.,3.,4.,5.,6.,7.,8.,9.,10.,11.,12.,13.,14.,15.,16.,17.,18.,19.,20.,21.,22.,23.;
	one_dim_rec_var=1,2,3,4,5,6,7,8,9,10;
	one_dim_rec_var_sng="Hello Wor";
	two_dim_rec_var_sng="abc",
				"bcd",
				"cde",
				"def",
				"efg",
				"fgh",
				"ghi",
				"hij",
				"jkl",
				"klm";
	char_var="z";
	rec_var_flt=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	rec_var_dbl=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	two_dim_rec_var=1.,2.0,3.,
			1.,2.1,3.,
			1.,2.2,3.,
			1.,2.3,3.,
			1.,2.4,3.,
			1.,2.5,3.,
			1.,2.6,3.,
			1.,2.7,3.,
			1.,2.8,3.,
			1.,2.9,3.;
	three_dim_rec_var= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				73,74,75,76,77,78,79,80;
	four_dim_rec_var= 	  1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12,
				 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24,
				 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36,
				 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48,
				 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60,
				 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72,
				 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84,
				 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96,
				 97, 98, 99,100,101,102,103,104,105,106,107,108,
				109,110,111,112,113,114,115,116,117,118,119,120,
				121,122,123,124,125,126,127,128,129,130,131,132,
				133,134,135,136,137,138,139,140,141,142,143,144,
				145,146,147,148,149,150,151,152,153,154,155,156,
				157,158,159,160,161,162,163,164,165,166,167,168,
				169,170,171,172,173,174,175,176,177,178,179,180,
				181,182,183,184,185,186,187,188,189,190,191,192,
				193,194,195,196,197,198,199,200,201,202,203,204,
				205,206,207,208,209,210,211,212,213,214,215,216,
				217,218,219,220,221,222,223,224,225,226,227,228,
				229,230,231,232,233,234,235,236,237,238,239,240;
}

