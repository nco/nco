// -*-C++-*-
// Purpose: CDL file to generate netCDF4 test file for vlen types

// Created: 20180413 based on buggy.cdl

// Usage:
// NB: ncgen arguments depend on version:
// "-k netCDF-4" for netCDF >= 3.6.3, "-k hdf5" for netCDF < 3.6.3
// "-k netCDF-4 classic model" for netCDF >= 3.6.3, "-k hdf5-nc3" for netCDF < 3.6.3
// ncgen -k netCDF-4 -b -o ~/nco/data/vlen.nc ~/nco/data/vlen.cdl
// scp ~/nco/data/vlen.cdl givre.ess.uci.edu:nco/data
// scp ~/nco/data/vlen.nc dust.ess.uci.edu:/var/www/html/nco
// scp dust.ess.uci.edu:/var/www/html/nco/vlen.nc ~/nco/data

netcdf vlen {

 types:
  int(*) vlen_int_t; // Declare "base-type" of vlen_int
  char(*) vlen_chr_t;
  string(*) vlen_sng_t; 
 dimensions:
  lat=2;

 variables:
  int one;
  
  vlen_int_t vlen_1D;
  vlen_1D:_FillValue={-999}; // vlen data MUST BE enclosed in braces
  vlen_int_t vlen_2D(lat);
  vlen_2D:_FillValue={-999};

  vlen_sng_t vlen_sng(lat);
 data:
  one=1;
  vlen_1D={17,18,19};
  vlen_2D={17,18,19},{1,2,3,4,5,6,7,_,9,_};
  vlen_sng={"one","two","three"},{"four,five"};

} // end root group
