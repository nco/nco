// Generate netCDF file with:
// ncgen -k netCDF-4 -b -o ~/nco/data/obs.nc ~/nco/data/obs.cdl

netcdf obs {
  dimensions:
  time=4;
  variables:
  float t(time);
  data:
  t=5,5,5,5;
 
} // end root group
