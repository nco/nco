netcdf snc_ncwa {

// global attributes:
		:institution = "NCAR (National Center for Atmospheric Research) Boulder, CO, USA" ;
		:institute_id = "NCAR" ;
		:experiment_id = "historical" ;
		:source = "CCSM4" ;
		:model_id = "CCSM4" ;
		:forcing = "Sl GHG Vl SS Ds SD BC MD OC Oz AA LU" ;
		:parent_experiment_id = "piControl" ;
		:parent_experiment_rip = "r1i1p1" ;
		:branch_time = 937. ;
		:contact = "cesm_data@ucar.edu" ;
		:references = "Gent P. R., et.al. 2011: The Community Climate System Model version 4. J. Climate, doi: 10.1175/2011JCLI4083.1" ;
		:initialization_method = 1 ;
		:physics_version = 1 ;
		:tracking_id = "a905e243-27f1-4172-93f0-820be7cbecf0" ;
		:acknowledgements = "The CESM project is supported by the National Science Foundation and the Office of Science (BER) of the U.S. Department of Energy. NCAR is sponsored by the National Science Foundation. Computing resources were provided by the Climate Simulation Laboratory at the NCAR Computational and Information Systems Laboratory (CISL), sponsored by the National Science Foundation and other agencies." ;
		:cesm_casename = "b40.20th.track1.1deg.008" ;
		:cesm_repotag = "ccsm4_0_beta43" ;
		:cesm_compset = "B20TRCN" ;
		:resolution = "f09_g16 (0.9x1.25_gx1v6)" ;
		:forcing_note = "Additional information on the external forcings used in this experiment can be found at http://www.cesm.ucar.edu/CMIP5/forcing_information" ;
		:processed_by = "strandwg on silver.cgd.ucar.edu at 20120406  -155645.062" ;
		:processing_code_information = "Last Changed Rev: 677 Last Changed Date: 2012-04-05 11:56:11 -0600 (Thu, 05 Apr 2012) Repository UUID: d2181dbe-5796-6825-dc7f-cbd98591f93d" ;
		:product = "output" ;
		:experiment = "historical" ;
		:frequency = "mon" ;
		:creation_date = "2012-04-06T21:56:48Z" ;
		:history = "Tue Aug 27 14:54:01 2013: ncecat --gag snc_LImon_CCSM4_historical_r1i1p1_199001-200512.nc snc_LImon_CESM1-BGC_esmHistorical_r1i1p1_199001-200512.nc snc_LImon_CESM1-BGC_historical_r1i1p1_199001-200512.nc snc_LImon_CESM1-CAM5_historical_r1i1p1_199001-200512.nc snc_LImon_CESM1-FASTCHEM_historical_r1i1p1_199001-200512.nc snc_LImon_CESM1-WACCM_historical_r1i1p1_199001-200512.nc snc.nc\nSun Dec 30 18:36:26 2012: ncks -d time,1990-01-01 00:00:0.0, /media/grele_data/wenshan/cesm/historical-exp/snc_LImon_CCSM4_historical_r1i1p1_185001-200512.nc /media/grele_data/wenshan/cesm/historical-exp/snc_LImon_CCSM4_historical_r1i1p1_199001-200512.nc\n2012-04-06T21:56:48Z CMOR rewrote data to comply with CF standards and CMIP5 requirements." ;
		:Conventions = "CF-1.4" ;
		:project_id = "CMIP5" ;
		:table_id = "Table LImon (12 January 2012) 429410275cb5466e41180ad9466db1bf" ;
		:title = "CCSM4 model output prepared for CMIP5 historical" ;
		:parent_experiment = "pre-industrial control" ;
		:modeling_realm = "landIce land" ;
		:realization = 1 ;
		:cmor_version = "2.8.1" ;
		:NCO = "20121231" ;
		:nco_openmp_thread_number = 1 ;

group: snc_LImon_CCSM4_historical_r1i1p1_199001-200512 {
  dimensions:
  	bnds = 2 ;
  	time = 192 ;
  variables:
  	double lat ;
  		lat:bounds = "lat_bnds" ;
  		lat:units = "degrees_north" ;
  		lat:axis = "Y" ;
  		lat:long_name = "latitude" ;
  		lat:standard_name = "latitude" ;
  	double lat_bnds(bnds) ;
  	double lon ;
  		lon:bounds = "lon_bnds" ;
  		lon:units = "degrees_east" ;
  		lon:axis = "X" ;
  		lon:long_name = "longitude" ;
  		lon:standard_name = "longitude" ;
  	double lon_bnds(bnds) ;
  	float snc(time) ;
  		snc:standard_name = "surface_snow_area_fraction" ;
  		snc:long_name = "Snow Area Fraction" ;
  		snc:comment = "FSNO, CMIP5_table_comment: Fraction of each grid cell that is occupied by snow that rests on land portion of cell." ;
  		snc:units = "%" ;
  		snc:original_name = "FSNO" ;
  		snc:cell_methods = "time: mean (interval: 30 days)" ;
  		snc:cell_measures = "area: areacella" ;
  		snc:history = "2012-04-06T21:56:45Z altered by CMOR: replaced missing value flag (1e+36) with standard missing value (1e+20)." ;
  		snc:missing_value = 1.e+20f ;
  		snc:_FillValue = 1.e+20f ;
  		snc:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_landIce_fx_CCSM4_historical_r0i0p0.nc areacella: areacella_fx_CCSM4_historical_r0i0p0.nc" ;
  	double time(time) ;
  		time:bounds = "time_bnds" ;
  		time:units = "days since 1850-01-01 00:00:00" ;
  		time:calendar = "noleap" ;
  		time:axis = "T" ;
  		time:long_name = "time" ;
  		time:standard_name = "time" ;
  	double time_bnds(time, bnds) ;

  // group attributes:
  		:institution = "NCAR (National Center for Atmospheric Research) Boulder, CO, USA" ;
  		:institute_id = "NCAR" ;
  		:experiment_id = "historical" ;
  		:source = "CCSM4" ;
  		:model_id = "CCSM4" ;
  		:forcing = "Sl GHG Vl SS Ds SD BC MD OC Oz AA LU" ;
  		:parent_experiment_id = "piControl" ;
  		:parent_experiment_rip = "r1i1p1" ;
  		:branch_time = 937. ;
  		:contact = "cesm_data@ucar.edu" ;
  		:references = "Gent P. R., et.al. 2011: The Community Climate System Model version 4. J. Climate, doi: 10.1175/2011JCLI4083.1" ;
  		:initialization_method = 1 ;
  		:physics_version = 1 ;
  		:tracking_id = "a905e243-27f1-4172-93f0-820be7cbecf0" ;
  		:acknowledgements = "The CESM project is supported by the National Science Foundation and the Office of Science (BER) of the U.S. Department of Energy. NCAR is sponsored by the National Science Foundation. Computing resources were provided by the Climate Simulation Laboratory at the NCAR Computational and Information Systems Laboratory (CISL), sponsored by the National Science Foundation and other agencies." ;
  		:cesm_casename = "b40.20th.track1.1deg.008" ;
  		:cesm_repotag = "ccsm4_0_beta43" ;
  		:cesm_compset = "B20TRCN" ;
  		:resolution = "f09_g16 (0.9x1.25_gx1v6)" ;
  		:forcing_note = "Additional information on the external forcings used in this experiment can be found at http://www.cesm.ucar.edu/CMIP5/forcing_information" ;
  		:processed_by = "strandwg on silver.cgd.ucar.edu at 20120406  -155645.062" ;
  		:processing_code_information = "Last Changed Rev: 677 Last Changed Date: 2012-04-05 11:56:11 -0600 (Thu, 05 Apr 2012) Repository UUID: d2181dbe-5796-6825-dc7f-cbd98591f93d" ;
  		:product = "output" ;
  		:experiment = "historical" ;
  		:frequency = "mon" ;
  		:creation_date = "2012-04-06T21:56:48Z" ;
  		:history = "Sun Dec 30 18:36:26 2012: ncks -d time,1990-01-01 00:00:0.0, /media/grele_data/wenshan/cesm/historical-exp/snc_LImon_CCSM4_historical_r1i1p1_185001-200512.nc /media/grele_data/wenshan/cesm/historical-exp/snc_LImon_CCSM4_historical_r1i1p1_199001-200512.nc\n2012-04-06T21:56:48Z CMOR rewrote data to comply with CF standards and CMIP5 requirements." ;
  		:Conventions = "CF-1.4" ;
  		:project_id = "CMIP5" ;
  		:table_id = "Table LImon (12 January 2012) 429410275cb5466e41180ad9466db1bf" ;
  		:title = "CCSM4 model output prepared for CMIP5 historical" ;
  		:parent_experiment = "pre-industrial control" ;
  		:modeling_realm = "landIce land" ;
  		:realization = 1 ;
  		:cmor_version = "2.8.1" ;
  		:NCO = "20121231" ;
  data:

   lat = 0 ;

   lat_bnds = -0.46875, 0.46875 ;

   lon = 179.375 ;

   lon_bnds = 178.752170138889, 180 ;

   snc = 61.37692, 60.05015, 58.4291, 52.22442, 45.59546, 38.34413, 33.19439, 
      32.58879, 36.96843, 46.77308, 55.4712, 60.32861, 61.04955, 60.44368, 
      57.63164, 52.03623, 44.6402, 37.95646, 33.34058, 32.47639, 35.50756, 
      46.31984, 53.72991, 58.95955, 60.95681, 61.11084, 57.52742, 51.32803, 
      45.14587, 40.29467, 33.73788, 32.70026, 37.01862, 45.55758, 54.71373, 
      59.162, 60.49402, 60.44479, 58.98337, 52.96589, 45.39301, 38.34033, 
      33.43645, 33.21604, 36.51387, 46.52538, 54.32355, 58.58232, 60.87978, 
      61.41938, 57.53942, 51.85412, 45.21275, 39.17278, 34.27933, 33.29999, 
      38.14444, 45.14943, 53.41065, 59.09114, 60.27861, 59.60844, 56.82986, 
      51.97681, 45.15635, 39.0167, 33.56191, 32.95903, 37.38646, 46.47746, 
      55.41323, 58.8252, 60.78623, 60.38117, 57.39877, 51.70517, 45.06911, 
      38.33918, 33.48069, 32.87983, 35.75778, 45.74866, 54.30301, 59.07576, 
      61.49643, 60.46125, 58.06967, 52.55259, 45.21442, 38.55085, 33.19324, 
      32.48174, 36.98698, 45.74392, 54.11422, 59.98495, 61.07553, 60.54321, 
      57.67136, 52.29048, 45.42659, 38.75619, 34.01928, 33.5902, 36.57975, 
      46.28279, 53.94093, 59.1823, 59.90117, 60.60514, 58.14232, 51.95426, 
      45.31351, 38.22518, 33.69085, 32.81738, 36.91416, 45.93295, 53.72042, 
      58.92241, 60.5704, 59.9584, 57.54922, 51.54271, 44.41114, 37.51797, 
      33.28756, 32.99597, 34.97438, 43.05939, 53.61963, 58.91531, 60.3945, 
      61.40278, 57.09048, 48.77563, 43.52256, 36.93203, 33.11032, 32.41613, 
      35.42476, 46.7383, 54.30549, 59.32918, 61.34241, 60.01548, 57.78593, 
      51.88309, 44.22643, 36.99844, 32.54312, 32.08076, 35.33289, 43.7334, 
      52.8833, 59.13483, 60.68259, 59.88637, 56.71269, 50.60006, 44.79, 
      38.0248, 32.8781, 32.3756, 36.24483, 44.34415, 54.8398, 59.24604, 
      60.13624, 60.5146, 57.35886, 51.2986, 44.53012, 38.94698, 32.69814, 
      32.66948, 36.62969, 45.27304, 53.99754, 57.90419, 61.03916, 59.86766, 
      55.66969, 51.11906, 44.3401, 38.34132, 33.50579, 32.66288, 36.10672, 
      46.07471, 53.37682, 59.08301 ;

   time = 51115.5, 51145, 51174.5, 51205, 51235.5, 51266, 51296.5, 51327.5, 
      51358, 51388.5, 51419, 51449.5, 51480.5, 51510, 51539.5, 51570, 
      51600.5, 51631, 51661.5, 51692.5, 51723, 51753.5, 51784, 51814.5, 
      51845.5, 51875, 51904.5, 51935, 51965.5, 51996, 52026.5, 52057.5, 
      52088, 52118.5, 52149, 52179.5, 52210.5, 52240, 52269.5, 52300, 
      52330.5, 52361, 52391.5, 52422.5, 52453, 52483.5, 52514, 52544.5, 
      52575.5, 52605, 52634.5, 52665, 52695.5, 52726, 52756.5, 52787.5, 
      52818, 52848.5, 52879, 52909.5, 52940.5, 52970, 52999.5, 53030, 
      53060.5, 53091, 53121.5, 53152.5, 53183, 53213.5, 53244, 53274.5, 
      53305.5, 53335, 53364.5, 53395, 53425.5, 53456, 53486.5, 53517.5, 
      53548, 53578.5, 53609, 53639.5, 53670.5, 53700, 53729.5, 53760, 
      53790.5, 53821, 53851.5, 53882.5, 53913, 53943.5, 53974, 54004.5, 
      54035.5, 54065, 54094.5, 54125, 54155.5, 54186, 54216.5, 54247.5, 
      54278, 54308.5, 54339, 54369.5, 54400.5, 54430, 54459.5, 54490, 
      54520.5, 54551, 54581.5, 54612.5, 54643, 54673.5, 54704, 54734.5, 
      54765.5, 54795, 54824.5, 54855, 54885.5, 54916, 54946.5, 54977.5, 
      55008, 55038.5, 55069, 55099.5, 55130.5, 55160, 55189.5, 55220, 
      55250.5, 55281, 55311.5, 55342.5, 55373, 55403.5, 55434, 55464.5, 
      55495.5, 55525, 55554.5, 55585, 55615.5, 55646, 55676.5, 55707.5, 
      55738, 55768.5, 55799, 55829.5, 55860.5, 55890, 55919.5, 55950, 
      55980.5, 56011, 56041.5, 56072.5, 56103, 56133.5, 56164, 56194.5, 
      56225.5, 56255, 56284.5, 56315, 56345.5, 56376, 56406.5, 56437.5, 
      56468, 56498.5, 56529, 56559.5, 56590.5, 56620, 56649.5, 56680, 
      56710.5, 56741, 56771.5, 56802.5, 56833, 56863.5, 56894, 56924.5 ;

   time_bnds =
  51100, 51131,
  51131, 51159,
  51159, 51190,
  51190, 51220,
  51220, 51251,
  51251, 51281,
  51281, 51312,
  51312, 51343,
  51343, 51373,
  51373, 51404,
  51404, 51434,
  51434, 51465,
  51465, 51496,
  51496, 51524,
  51524, 51555,
  51555, 51585,
  51585, 51616,
  51616, 51646,
  51646, 51677,
  51677, 51708,
  51708, 51738,
  51738, 51769,
  51769, 51799,
  51799, 51830,
  51830, 51861,
  51861, 51889,
  51889, 51920,
  51920, 51950,
  51950, 51981,
  51981, 52011,
  52011, 52042,
  52042, 52073,
  52073, 52103,
  52103, 52134,
  52134, 52164,
  52164, 52195,
  52195, 52226,
  52226, 52254,
  52254, 52285,
  52285, 52315,
  52315, 52346,
  52346, 52376,
  52376, 52407,
  52407, 52438,
  52438, 52468,
  52468, 52499,
  52499, 52529,
  52529, 52560,
  52560, 52591,
  52591, 52619,
  52619, 52650,
  52650, 52680,
  52680, 52711,
  52711, 52741,
  52741, 52772,
  52772, 52803,
  52803, 52833,
  52833, 52864,
  52864, 52894,
  52894, 52925,
  52925, 52956,
  52956, 52984,
  52984, 53015,
  53015, 53045,
  53045, 53076,
  53076, 53106,
  53106, 53137,
  53137, 53168,
  53168, 53198,
  53198, 53229,
  53229, 53259,
  53259, 53290,
  53290, 53321,
  53321, 53349,
  53349, 53380,
  53380, 53410,
  53410, 53441,
  53441, 53471,
  53471, 53502,
  53502, 53533,
  53533, 53563,
  53563, 53594,
  53594, 53624,
  53624, 53655,
  53655, 53686,
  53686, 53714,
  53714, 53745,
  53745, 53775,
  53775, 53806,
  53806, 53836,
  53836, 53867,
  53867, 53898,
  53898, 53928,
  53928, 53959,
  53959, 53989,
  53989, 54020,
  54020, 54051,
  54051, 54079,
  54079, 54110,
  54110, 54140,
  54140, 54171,
  54171, 54201,
  54201, 54232,
  54232, 54263,
  54263, 54293,
  54293, 54324,
  54324, 54354,
  54354, 54385,
  54385, 54416,
  54416, 54444,
  54444, 54475,
  54475, 54505,
  54505, 54536,
  54536, 54566,
  54566, 54597,
  54597, 54628,
  54628, 54658,
  54658, 54689,
  54689, 54719,
  54719, 54750,
  54750, 54781,
  54781, 54809,
  54809, 54840,
  54840, 54870,
  54870, 54901,
  54901, 54931,
  54931, 54962,
  54962, 54993,
  54993, 55023,
  55023, 55054,
  55054, 55084,
  55084, 55115,
  55115, 55146,
  55146, 55174,
  55174, 55205,
  55205, 55235,
  55235, 55266,
  55266, 55296,
  55296, 55327,
  55327, 55358,
  55358, 55388,
  55388, 55419,
  55419, 55449,
  55449, 55480,
  55480, 55511,
  55511, 55539,
  55539, 55570,
  55570, 55600,
  55600, 55631,
  55631, 55661,
  55661, 55692,
  55692, 55723,
  55723, 55753,
  55753, 55784,
  55784, 55814,
  55814, 55845,
  55845, 55876,
  55876, 55904,
  55904, 55935,
  55935, 55965,
  55965, 55996,
  55996, 56026,
  56026, 56057,
  56057, 56088,
  56088, 56118,
  56118, 56149,
  56149, 56179,
  56179, 56210,
  56210, 56241,
  56241, 56269,
  56269, 56300,
  56300, 56330,
  56330, 56361,
  56361, 56391,
  56391, 56422,
  56422, 56453,
  56453, 56483,
  56483, 56514,
  56514, 56544,
  56544, 56575,
  56575, 56606,
  56606, 56634,
  56634, 56665,
  56665, 56695,
  56695, 56726,
  56726, 56756,
  56756, 56787,
  56787, 56818,
  56818, 56848,
  56848, 56879,
  56879, 56909,
  56909, 56940 ;
  } // group snc_LImon_CCSM4_historical_r1i1p1_199001-200512

group: snc_LImon_CESM1-BGC_esmHistorical_r1i1p1_199001-200512 {
  dimensions:
  	bnds = 2 ;
  	time = 192 ;
  variables:
  	double lat ;
  		lat:bounds = "lat_bnds" ;
  		lat:units = "degrees_north" ;
  		lat:axis = "Y" ;
  		lat:long_name = "latitude" ;
  		lat:standard_name = "latitude" ;
  	double lat_bnds(bnds) ;
  	double lon ;
  		lon:bounds = "lon_bnds" ;
  		lon:units = "degrees_east" ;
  		lon:axis = "X" ;
  		lon:long_name = "longitude" ;
  		lon:standard_name = "longitude" ;
  	double lon_bnds(bnds) ;
  	float snc(time) ;
  		snc:standard_name = "surface_snow_area_fraction" ;
  		snc:long_name = "Snow Area Fraction" ;
  		snc:comment = "FSNO, CMIP5_table_comment: Fraction of each grid cell that is occupied by snow that rests on land portion of cell." ;
  		snc:units = "%" ;
  		snc:original_name = "FSNO" ;
  		snc:cell_methods = "time: mean (interval: 30 days)" ;
  		snc:cell_measures = "area: areacella" ;
  		snc:history = "2012-05-09T19:56:59Z altered by CMOR: replaced missing value flag (1e+36) with standard missing value (1e+20)." ;
  		snc:missing_value = 1.e+20f ;
  		snc:_FillValue = 1.e+20f ;
  		snc:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_landIce_fx_CESM1-BGC_esmHistorical_r0i0p0.nc areacella: areacella_fx_CESM1-BGC_esmHistorical_r0i0p0.nc" ;
  	double time(time) ;
  		time:bounds = "time_bnds" ;
  		time:units = "days since 1850-01-01 00:00:00" ;
  		time:calendar = "noleap" ;
  		time:axis = "T" ;
  		time:long_name = "time" ;
  		time:standard_name = "time" ;
  	double time_bnds(time, bnds) ;

  // group attributes:
  		:institution = "NSF/DOE NCAR (National Center for Atmospheric Research) Boulder, CO, USA" ;
  		:institute_id = "NSF-DOE-NCAR" ;
  		:experiment_id = "esmHistorical" ;
  		:source = "CESM1-BGC" ;
  		:model_id = "CESM1-BGC" ;
  		:forcing = "Sl GHG Vl SS Ds SD BC MD OC Oz AA LU" ;
  		:parent_experiment_id = "piControl" ;
  		:parent_experiment_rip = "r1i1p1" ;
  		:branch_time = 1. ;
  		:contact = "cesm_data@ucar.edu" ;
  		:comment = "CESM home page: http://www.cesm.ucar.edu" ;
  		:references = "TBD\n See also http://www.cesm.ucar.edu/publications" ;
  		:initialization_method = 1 ;
  		:physics_version = 1 ;
  		:tracking_id = "c763c1db-4d63-4268-aa34-b1a9ca11cb75" ;
  		:acknowledgements = "The CESM project is supported by the National Science Foundation and the Office of Science (BER) of the U.S. Department of Energy. NCAR is sponsored by the National Science Foundation. Computing resources were provided by the Climate Simulation Laboratory at the NCAR Computational and Information Systems Laboratory (CISL), sponsored by the National Science Foundation and other agencies." ;
  		:cesm_casename = "b40.20th.1deg.coup.001" ;
  		:cesm_repotag = "unknown" ;
  		:cesm_compset = "unknown" ;
  		:resolution = "f09_g16 (0.9x1.25_gx1v6)" ;
  		:forcing_note = "Additional information on the external forcings used in this experiment can be found at http://www.cesm.ucar.edu/CMIP5/forcing_information" ;
  		:processed_by = "strandwg on silver.cgd.ucar.edu at 20120509  -135659.177" ;
  		:processing_code_information = "Last Changed Rev: 757 Last Changed Date: 2012-05-09 13:01:12 -0600 (Wed, 09 May 2012) Repository UUID: d2181dbe-5796-6825-dc7f-cbd98591f93d" ;
  		:product = "output" ;
  		:experiment = "ESM historical" ;
  		:frequency = "mon" ;
  		:creation_date = "2012-05-09T19:57:12Z" ;
  		:history = "Sun Dec 30 18:37:17 2012: ncks -d time,1990-01-01 00:00:0.0, /media/grele_data/wenshan/cesm/historical-exp/snc_LImon_CESM1-BGC_esmHistorical_r1i1p1_185001-200512.nc /media/grele_data/wenshan/cesm/historical-exp/snc_LImon_CESM1-BGC_esmHistorical_r1i1p1_199001-200512.nc\n2012-05-09T19:57:12Z CMOR rewrote data to comply with CF standards and CMIP5 requirements." ;
  		:Conventions = "CF-1.4" ;
  		:project_id = "CMIP5" ;
  		:table_id = "Table LImon (12 January 2012) 429410275cb5466e41180ad9466db1bf" ;
  		:title = "CESM1-BGC model output prepared for CMIP5 ESM historical" ;
  		:parent_experiment = "pre-industrial control" ;
  		:modeling_realm = "landIce land" ;
  		:realization = 1 ;
  		:cmor_version = "2.8.1" ;
  		:NCO = "20121231" ;
  data:

   lat = 0 ;

   lat_bnds = -0.46875, 0.46875 ;

   lon = 179.375 ;

   lon_bnds = 178.752170138889, 180 ;

   snc = 60.42937, 60.64738, 57.30071, 51.4353, 45.43332, 39.52806, 34.66951, 
      33.13662, 36.25096, 46.04024, 53.33717, 59.30924, 60.99267, 59.43881, 
      57.94574, 51.67841, 44.91564, 39.39613, 34.42404, 33.53218, 36.72351, 
      47.10626, 54.4623, 58.49553, 59.56153, 59.97334, 57.89266, 52.57605, 
      45.66745, 38.9083, 34.23455, 34.08851, 38.44006, 47.2091, 55.48892, 
      60.75134, 61.30203, 61.29112, 60.0729, 54.08234, 46.12404, 38.92447, 
      34.04529, 33.68865, 37.31947, 45.64073, 55.82588, 60.10115, 61.4198, 
      59.77499, 56.8927, 51.5806, 45.45844, 38.9374, 34.54553, 33.49256, 
      36.34779, 46.30656, 53.9354, 58.88356, 60.45415, 60.14672, 57.57286, 
      52.50472, 46.36785, 39.8609, 33.63399, 33.20422, 35.44655, 44.78173, 
      53.92061, 59.74142, 60.50524, 60.10552, 58.04763, 51.95174, 45.57401, 
      39.92517, 34.07393, 33.18673, 36.03875, 46.52081, 54.78568, 59.38622, 
      60.48057, 59.2347, 56.71712, 52.24715, 46.07843, 38.27985, 33.38749, 
      33.0439, 35.73171, 45.55057, 53.66148, 58.66822, 61.14587, 61.68203, 
      57.431, 50.35966, 44.36692, 38.19395, 33.53297, 33.26769, 35.39089, 
      45.34281, 54.08255, 59.35721, 61.94003, 60.47675, 56.81584, 51.78187, 
      45.66067, 39.36295, 33.72239, 33.26345, 36.18309, 44.39331, 52.50751, 
      59.50554, 61.95173, 60.64665, 57.34688, 51.2981, 45.21524, 38.18364, 
      33.42353, 32.79172, 35.11573, 43.63971, 53.21791, 58.21271, 59.6288, 
      61.27858, 56.47172, 50.35821, 43.80642, 37.97486, 33.80445, 33.41068, 
      35.89848, 46.58085, 54.50834, 59.01017, 61.5377, 60.76017, 57.91518, 
      51.82125, 43.89352, 38.06473, 33.38121, 32.91643, 35.2864, 45.38606, 
      53.46272, 59.2138, 60.37124, 59.06458, 55.75334, 50.40107, 44.48877, 
      38.5047, 33.78501, 33.20532, 36.02801, 43.41591, 53.39999, 58.97802, 
      60.57231, 59.36517, 55.10088, 49.68346, 44.11604, 38.80204, 33.5981, 
      32.79944, 36.32286, 44.73896, 53.55066, 58.98016, 60.80568, 59.11828, 
      55.20478, 50.08527, 44.43622, 38.27273, 33.41451, 32.98672, 35.45163, 
      44.04631, 52.83684, 59.77518 ;

   time = 51115.5, 51145, 51174.5, 51205, 51235.5, 51266, 51296.5, 51327.5, 
      51358, 51388.5, 51419, 51449.5, 51480.5, 51510, 51539.5, 51570, 
      51600.5, 51631, 51661.5, 51692.5, 51723, 51753.5, 51784, 51814.5, 
      51845.5, 51875, 51904.5, 51935, 51965.5, 51996, 52026.5, 52057.5, 
      52088, 52118.5, 52149, 52179.5, 52210.5, 52240, 52269.5, 52300, 
      52330.5, 52361, 52391.5, 52422.5, 52453, 52483.5, 52514, 52544.5, 
      52575.5, 52605, 52634.5, 52665, 52695.5, 52726, 52756.5, 52787.5, 
      52818, 52848.5, 52879, 52909.5, 52940.5, 52970, 52999.5, 53030, 
      53060.5, 53091, 53121.5, 53152.5, 53183, 53213.5, 53244, 53274.5, 
      53305.5, 53335, 53364.5, 53395, 53425.5, 53456, 53486.5, 53517.5, 
      53548, 53578.5, 53609, 53639.5, 53670.5, 53700, 53729.5, 53760, 
      53790.5, 53821, 53851.5, 53882.5, 53913, 53943.5, 53974, 54004.5, 
      54035.5, 54065, 54094.5, 54125, 54155.5, 54186, 54216.5, 54247.5, 
      54278, 54308.5, 54339, 54369.5, 54400.5, 54430, 54459.5, 54490, 
      54520.5, 54551, 54581.5, 54612.5, 54643, 54673.5, 54704, 54734.5, 
      54765.5, 54795, 54824.5, 54855, 54885.5, 54916, 54946.5, 54977.5, 
      55008, 55038.5, 55069, 55099.5, 55130.5, 55160, 55189.5, 55220, 
      55250.5, 55281, 55311.5, 55342.5, 55373, 55403.5, 55434, 55464.5, 
      55495.5, 55525, 55554.5, 55585, 55615.5, 55646, 55676.5, 55707.5, 
      55738, 55768.5, 55799, 55829.5, 55860.5, 55890, 55919.5, 55950, 
      55980.5, 56011, 56041.5, 56072.5, 56103, 56133.5, 56164, 56194.5, 
      56225.5, 56255, 56284.5, 56315, 56345.5, 56376, 56406.5, 56437.5, 
      56468, 56498.5, 56529, 56559.5, 56590.5, 56620, 56649.5, 56680, 
      56710.5, 56741, 56771.5, 56802.5, 56833, 56863.5, 56894, 56924.5 ;

   time_bnds =
  51100, 51131,
  51131, 51159,
  51159, 51190,
  51190, 51220,
  51220, 51251,
  51251, 51281,
  51281, 51312,
  51312, 51343,
  51343, 51373,
  51373, 51404,
  51404, 51434,
  51434, 51465,
  51465, 51496,
  51496, 51524,
  51524, 51555,
  51555, 51585,
  51585, 51616,
  51616, 51646,
  51646, 51677,
  51677, 51708,
  51708, 51738,
  51738, 51769,
  51769, 51799,
  51799, 51830,
  51830, 51861,
  51861, 51889,
  51889, 51920,
  51920, 51950,
  51950, 51981,
  51981, 52011,
  52011, 52042,
  52042, 52073,
  52073, 52103,
  52103, 52134,
  52134, 52164,
  52164, 52195,
  52195, 52226,
  52226, 52254,
  52254, 52285,
  52285, 52315,
  52315, 52346,
  52346, 52376,
  52376, 52407,
  52407, 52438,
  52438, 52468,
  52468, 52499,
  52499, 52529,
  52529, 52560,
  52560, 52591,
  52591, 52619,
  52619, 52650,
  52650, 52680,
  52680, 52711,
  52711, 52741,
  52741, 52772,
  52772, 52803,
  52803, 52833,
  52833, 52864,
  52864, 52894,
  52894, 52925,
  52925, 52956,
  52956, 52984,
  52984, 53015,
  53015, 53045,
  53045, 53076,
  53076, 53106,
  53106, 53137,
  53137, 53168,
  53168, 53198,
  53198, 53229,
  53229, 53259,
  53259, 53290,
  53290, 53321,
  53321, 53349,
  53349, 53380,
  53380, 53410,
  53410, 53441,
  53441, 53471,
  53471, 53502,
  53502, 53533,
  53533, 53563,
  53563, 53594,
  53594, 53624,
  53624, 53655,
  53655, 53686,
  53686, 53714,
  53714, 53745,
  53745, 53775,
  53775, 53806,
  53806, 53836,
  53836, 53867,
  53867, 53898,
  53898, 53928,
  53928, 53959,
  53959, 53989,
  53989, 54020,
  54020, 54051,
  54051, 54079,
  54079, 54110,
  54110, 54140,
  54140, 54171,
  54171, 54201,
  54201, 54232,
  54232, 54263,
  54263, 54293,
  54293, 54324,
  54324, 54354,
  54354, 54385,
  54385, 54416,
  54416, 54444,
  54444, 54475,
  54475, 54505,
  54505, 54536,
  54536, 54566,
  54566, 54597,
  54597, 54628,
  54628, 54658,
  54658, 54689,
  54689, 54719,
  54719, 54750,
  54750, 54781,
  54781, 54809,
  54809, 54840,
  54840, 54870,
  54870, 54901,
  54901, 54931,
  54931, 54962,
  54962, 54993,
  54993, 55023,
  55023, 55054,
  55054, 55084,
  55084, 55115,
  55115, 55146,
  55146, 55174,
  55174, 55205,
  55205, 55235,
  55235, 55266,
  55266, 55296,
  55296, 55327,
  55327, 55358,
  55358, 55388,
  55388, 55419,
  55419, 55449,
  55449, 55480,
  55480, 55511,
  55511, 55539,
  55539, 55570,
  55570, 55600,
  55600, 55631,
  55631, 55661,
  55661, 55692,
  55692, 55723,
  55723, 55753,
  55753, 55784,
  55784, 55814,
  55814, 55845,
  55845, 55876,
  55876, 55904,
  55904, 55935,
  55935, 55965,
  55965, 55996,
  55996, 56026,
  56026, 56057,
  56057, 56088,
  56088, 56118,
  56118, 56149,
  56149, 56179,
  56179, 56210,
  56210, 56241,
  56241, 56269,
  56269, 56300,
  56300, 56330,
  56330, 56361,
  56361, 56391,
  56391, 56422,
  56422, 56453,
  56453, 56483,
  56483, 56514,
  56514, 56544,
  56544, 56575,
  56575, 56606,
  56606, 56634,
  56634, 56665,
  56665, 56695,
  56695, 56726,
  56726, 56756,
  56756, 56787,
  56787, 56818,
  56818, 56848,
  56848, 56879,
  56879, 56909,
  56909, 56940 ;
  } // group snc_LImon_CESM1-BGC_esmHistorical_r1i1p1_199001-200512

group: snc_LImon_CESM1-BGC_historical_r1i1p1_199001-200512 {
  dimensions:
  	bnds = 2 ;
  	time = 192 ;
  variables:
  	double lat ;
  		lat:bounds = "lat_bnds" ;
  		lat:units = "degrees_north" ;
  		lat:axis = "Y" ;
  		lat:long_name = "latitude" ;
  		lat:standard_name = "latitude" ;
  	double lat_bnds(bnds) ;
  	double lon ;
  		lon:bounds = "lon_bnds" ;
  		lon:units = "degrees_east" ;
  		lon:axis = "X" ;
  		lon:long_name = "longitude" ;
  		lon:standard_name = "longitude" ;
  	double lon_bnds(bnds) ;
  	float snc(time) ;
  		snc:standard_name = "surface_snow_area_fraction" ;
  		snc:long_name = "Snow Area Fraction" ;
  		snc:comment = "FSNO, CMIP5_table_comment: Fraction of each grid cell that is occupied by snow that rests on land portion of cell." ;
  		snc:units = "%" ;
  		snc:original_name = "FSNO" ;
  		snc:cell_methods = "time: mean (interval: 30 days)" ;
  		snc:cell_measures = "area: areacella" ;
  		snc:history = "2012-05-09T19:57:50Z altered by CMOR: replaced missing value flag (1e+36) with standard missing value (1e+20)." ;
  		snc:missing_value = 1.e+20f ;
  		snc:_FillValue = 1.e+20f ;
  		snc:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_landIce_fx_CESM1-BGC_historical_r0i0p0.nc areacella: areacella_fx_CESM1-BGC_historical_r0i0p0.nc" ;
  	double time(time) ;
  		time:bounds = "time_bnds" ;
  		time:units = "days since 1850-01-01 00:00:00" ;
  		time:calendar = "noleap" ;
  		time:axis = "T" ;
  		time:long_name = "time" ;
  		time:standard_name = "time" ;
  	double time_bnds(time, bnds) ;

  // group attributes:
  		:institution = "NSF/DOE NCAR (National Center for Atmospheric Research) Boulder, CO, USA" ;
  		:institute_id = "NSF-DOE-NCAR" ;
  		:experiment_id = "historical" ;
  		:source = "CESM1-BGC" ;
  		:model_id = "CESM1-BGC" ;
  		:forcing = "Sl GHG Vl SS Ds SD BC MD OC Oz AA LU" ;
  		:parent_experiment_id = "piControl" ;
  		:parent_experiment_rip = "r1i1p1" ;
  		:branch_time = 1. ;
  		:contact = "cesm_data@ucar.edu" ;
  		:comment = "CESM home page: http://www.cesm.ucar.edu" ;
  		:references = "TBD\n See also http://www.cesm.ucar.edu/publications" ;
  		:initialization_method = 1 ;
  		:physics_version = 1 ;
  		:tracking_id = "1b9bc30c-5957-4e3f-999f-0a28b5f60139" ;
  		:acknowledgements = "The CESM project is supported by the National Science Foundation and the Office of Science (BER) of the U.S. Department of Energy. NCAR is sponsored by the National Science Foundation. Computing resources were provided by the Climate Simulation Laboratory at the NCAR Computational and Information Systems Laboratory (CISL), sponsored by the National Science Foundation and other agencies." ;
  		:cesm_casename = "b40.20th.1deg.bdrd.001" ;
  		:cesm_repotag = "unknown" ;
  		:cesm_compset = "unknown" ;
  		:resolution = "f09_g16 (0.9x1.25_gx1v6)" ;
  		:forcing_note = "Additional information on the external forcings used in this experiment can be found at http://www.cesm.ucar.edu/CMIP5/forcing_information" ;
  		:processed_by = "strandwg on silver.cgd.ucar.edu at 20120509  -135750.546" ;
  		:processing_code_information = "Last Changed Rev: 757 Last Changed Date: 2012-05-09 13:01:12 -0600 (Wed, 09 May 2012) Repository UUID: d2181dbe-5796-6825-dc7f-cbd98591f93d" ;
  		:product = "output" ;
  		:experiment = "historical" ;
  		:frequency = "mon" ;
  		:creation_date = "2012-05-09T19:58:05Z" ;
  		:history = "Thu Jan 24 16:59:20 2013: ncks -d time,1990-01-01 00:00:0.0, snc_LImon_CESM1-BGC_historical_r1i1p1_185001-200512.nc snc_LImon_CESM1-BGC_historical_r1i1p1_199001-200512.nc\n2012-05-09T19:58:05Z CMOR rewrote data to comply with CF standards and CMIP5 requirements." ;
  		:Conventions = "CF-1.4" ;
  		:project_id = "CMIP5" ;
  		:table_id = "Table LImon (12 January 2012) 429410275cb5466e41180ad9466db1bf" ;
  		:title = "CESM1-BGC model output prepared for CMIP5 historical" ;
  		:parent_experiment = "pre-industrial control" ;
  		:modeling_realm = "landIce land" ;
  		:realization = 1 ;
  		:cmor_version = "2.8.1" ;
  		:NCO = "20130125" ;
  data:

   lat = 0 ;

   lat_bnds = -0.46875, 0.46875 ;

   lon = 179.375 ;

   lon_bnds = 178.752170138889, 180 ;

   snc = 60.81151, 60.83581, 57.40618, 50.77258, 45.05299, 38.55186, 
      33.70737, 33.04415, 35.72379, 47.15994, 53.97527, 58.59232, 62.0451, 
      60.02757, 57.57421, 52.67574, 45.38245, 38.96038, 33.7025, 33.30761, 
      36.09553, 45.33242, 53.43705, 59.69139, 60.2207, 59.44222, 57.08393, 
      51.60577, 45.91001, 40.35986, 35.51391, 33.55119, 37.95975, 46.05239, 
      55.25557, 60.17647, 61.67732, 61.58868, 57.89724, 51.44344, 45.45924, 
      39.27931, 33.92011, 33.49309, 37.62573, 45.77045, 54.64713, 60.00785, 
      62.98378, 60.98982, 57.44807, 53.21042, 45.43661, 38.67152, 33.94413, 
      33.15783, 35.94777, 44.61528, 54.27599, 58.80817, 61.2307, 59.79439, 
      57.08263, 50.52497, 44.07899, 38.27042, 33.51943, 32.94697, 35.40871, 
      45.28115, 53.79686, 59.03689, 60.84576, 59.65984, 57.90582, 52.30964, 
      45.07834, 39.25048, 33.8819, 33.14655, 35.57959, 44.89124, 54.50274, 
      58.59656, 60.65822, 59.59388, 56.29368, 50.73042, 43.93979, 37.35862, 
      33.44497, 32.98347, 36.43193, 44.7622, 54.04124, 58.71893, 59.85044, 
      60.0969, 57.5133, 51.66403, 45.28492, 38.6044, 34.07675, 33.54704, 
      36.35543, 43.59683, 52.81324, 59.19917, 62.49909, 59.65298, 55.79979, 
      51.49189, 46.20795, 39.5049, 34.17224, 33.11736, 37.46117, 44.75187, 
      53.72094, 59.15183, 61.0971, 59.81115, 56.52975, 51.89294, 45.86815, 
      38.33873, 33.06678, 32.81318, 35.49161, 45.98712, 53.63966, 59.74233, 
      61.00092, 61.10449, 57.47633, 51.74292, 45.13937, 37.65129, 33.35644, 
      33.50973, 35.10047, 44.06165, 54.06438, 60.30418, 61.70724, 61.21657, 
      58.94371, 52.51987, 45.48262, 38.52264, 33.92553, 32.91373, 35.71524, 
      46.23709, 53.22155, 58.81511, 59.43888, 59.1026, 56.43563, 50.23117, 
      43.67832, 37.89594, 33.47663, 32.65866, 35.80147, 45.50639, 52.66769, 
      58.6243, 60.40725, 59.98502, 57.12119, 51.65089, 45.57036, 38.15372, 
      32.98792, 32.49368, 35.69475, 45.33248, 52.4259, 57.92989, 60.0364, 
      59.07898, 56.09073, 50.74621, 43.55686, 37.64441, 33.23428, 32.99554, 
      36.66736, 44.9342, 54.54264, 58.61319 ;

   time = 51115.5, 51145, 51174.5, 51205, 51235.5, 51266, 51296.5, 51327.5, 
      51358, 51388.5, 51419, 51449.5, 51480.5, 51510, 51539.5, 51570, 
      51600.5, 51631, 51661.5, 51692.5, 51723, 51753.5, 51784, 51814.5, 
      51845.5, 51875, 51904.5, 51935, 51965.5, 51996, 52026.5, 52057.5, 
      52088, 52118.5, 52149, 52179.5, 52210.5, 52240, 52269.5, 52300, 
      52330.5, 52361, 52391.5, 52422.5, 52453, 52483.5, 52514, 52544.5, 
      52575.5, 52605, 52634.5, 52665, 52695.5, 52726, 52756.5, 52787.5, 
      52818, 52848.5, 52879, 52909.5, 52940.5, 52970, 52999.5, 53030, 
      53060.5, 53091, 53121.5, 53152.5, 53183, 53213.5, 53244, 53274.5, 
      53305.5, 53335, 53364.5, 53395, 53425.5, 53456, 53486.5, 53517.5, 
      53548, 53578.5, 53609, 53639.5, 53670.5, 53700, 53729.5, 53760, 
      53790.5, 53821, 53851.5, 53882.5, 53913, 53943.5, 53974, 54004.5, 
      54035.5, 54065, 54094.5, 54125, 54155.5, 54186, 54216.5, 54247.5, 
      54278, 54308.5, 54339, 54369.5, 54400.5, 54430, 54459.5, 54490, 
      54520.5, 54551, 54581.5, 54612.5, 54643, 54673.5, 54704, 54734.5, 
      54765.5, 54795, 54824.5, 54855, 54885.5, 54916, 54946.5, 54977.5, 
      55008, 55038.5, 55069, 55099.5, 55130.5, 55160, 55189.5, 55220, 
      55250.5, 55281, 55311.5, 55342.5, 55373, 55403.5, 55434, 55464.5, 
      55495.5, 55525, 55554.5, 55585, 55615.5, 55646, 55676.5, 55707.5, 
      55738, 55768.5, 55799, 55829.5, 55860.5, 55890, 55919.5, 55950, 
      55980.5, 56011, 56041.5, 56072.5, 56103, 56133.5, 56164, 56194.5, 
      56225.5, 56255, 56284.5, 56315, 56345.5, 56376, 56406.5, 56437.5, 
      56468, 56498.5, 56529, 56559.5, 56590.5, 56620, 56649.5, 56680, 
      56710.5, 56741, 56771.5, 56802.5, 56833, 56863.5, 56894, 56924.5 ;

   time_bnds =
  51100, 51131,
  51131, 51159,
  51159, 51190,
  51190, 51220,
  51220, 51251,
  51251, 51281,
  51281, 51312,
  51312, 51343,
  51343, 51373,
  51373, 51404,
  51404, 51434,
  51434, 51465,
  51465, 51496,
  51496, 51524,
  51524, 51555,
  51555, 51585,
  51585, 51616,
  51616, 51646,
  51646, 51677,
  51677, 51708,
  51708, 51738,
  51738, 51769,
  51769, 51799,
  51799, 51830,
  51830, 51861,
  51861, 51889,
  51889, 51920,
  51920, 51950,
  51950, 51981,
  51981, 52011,
  52011, 52042,
  52042, 52073,
  52073, 52103,
  52103, 52134,
  52134, 52164,
  52164, 52195,
  52195, 52226,
  52226, 52254,
  52254, 52285,
  52285, 52315,
  52315, 52346,
  52346, 52376,
  52376, 52407,
  52407, 52438,
  52438, 52468,
  52468, 52499,
  52499, 52529,
  52529, 52560,
  52560, 52591,
  52591, 52619,
  52619, 52650,
  52650, 52680,
  52680, 52711,
  52711, 52741,
  52741, 52772,
  52772, 52803,
  52803, 52833,
  52833, 52864,
  52864, 52894,
  52894, 52925,
  52925, 52956,
  52956, 52984,
  52984, 53015,
  53015, 53045,
  53045, 53076,
  53076, 53106,
  53106, 53137,
  53137, 53168,
  53168, 53198,
  53198, 53229,
  53229, 53259,
  53259, 53290,
  53290, 53321,
  53321, 53349,
  53349, 53380,
  53380, 53410,
  53410, 53441,
  53441, 53471,
  53471, 53502,
  53502, 53533,
  53533, 53563,
  53563, 53594,
  53594, 53624,
  53624, 53655,
  53655, 53686,
  53686, 53714,
  53714, 53745,
  53745, 53775,
  53775, 53806,
  53806, 53836,
  53836, 53867,
  53867, 53898,
  53898, 53928,
  53928, 53959,
  53959, 53989,
  53989, 54020,
  54020, 54051,
  54051, 54079,
  54079, 54110,
  54110, 54140,
  54140, 54171,
  54171, 54201,
  54201, 54232,
  54232, 54263,
  54263, 54293,
  54293, 54324,
  54324, 54354,
  54354, 54385,
  54385, 54416,
  54416, 54444,
  54444, 54475,
  54475, 54505,
  54505, 54536,
  54536, 54566,
  54566, 54597,
  54597, 54628,
  54628, 54658,
  54658, 54689,
  54689, 54719,
  54719, 54750,
  54750, 54781,
  54781, 54809,
  54809, 54840,
  54840, 54870,
  54870, 54901,
  54901, 54931,
  54931, 54962,
  54962, 54993,
  54993, 55023,
  55023, 55054,
  55054, 55084,
  55084, 55115,
  55115, 55146,
  55146, 55174,
  55174, 55205,
  55205, 55235,
  55235, 55266,
  55266, 55296,
  55296, 55327,
  55327, 55358,
  55358, 55388,
  55388, 55419,
  55419, 55449,
  55449, 55480,
  55480, 55511,
  55511, 55539,
  55539, 55570,
  55570, 55600,
  55600, 55631,
  55631, 55661,
  55661, 55692,
  55692, 55723,
  55723, 55753,
  55753, 55784,
  55784, 55814,
  55814, 55845,
  55845, 55876,
  55876, 55904,
  55904, 55935,
  55935, 55965,
  55965, 55996,
  55996, 56026,
  56026, 56057,
  56057, 56088,
  56088, 56118,
  56118, 56149,
  56149, 56179,
  56179, 56210,
  56210, 56241,
  56241, 56269,
  56269, 56300,
  56300, 56330,
  56330, 56361,
  56361, 56391,
  56391, 56422,
  56422, 56453,
  56453, 56483,
  56483, 56514,
  56514, 56544,
  56544, 56575,
  56575, 56606,
  56606, 56634,
  56634, 56665,
  56665, 56695,
  56695, 56726,
  56726, 56756,
  56756, 56787,
  56787, 56818,
  56818, 56848,
  56848, 56879,
  56879, 56909,
  56909, 56940 ;
  } // group snc_LImon_CESM1-BGC_historical_r1i1p1_199001-200512

group: snc_LImon_CESM1-CAM5_historical_r1i1p1_199001-200512 {
  dimensions:
  	bnds = 2 ;
  	time = 192 ;
  variables:
  	double lat ;
  		lat:bounds = "lat_bnds" ;
  		lat:units = "degrees_north" ;
  		lat:axis = "Y" ;
  		lat:long_name = "latitude" ;
  		lat:standard_name = "latitude" ;
  	double lat_bnds(bnds) ;
  	double lon ;
  		lon:bounds = "lon_bnds" ;
  		lon:units = "degrees_east" ;
  		lon:axis = "X" ;
  		lon:long_name = "longitude" ;
  		lon:standard_name = "longitude" ;
  	double lon_bnds(bnds) ;
  	float snc(time) ;
  		snc:standard_name = "surface_snow_area_fraction" ;
  		snc:long_name = "Snow Area Fraction" ;
  		snc:comment = "FSNO, CMIP5_table_comment: Fraction of each grid cell that is occupied by snow that rests on land portion of cell." ;
  		snc:units = "%" ;
  		snc:original_name = "FSNO" ;
  		snc:cell_methods = "time: mean (interval: 30 days)" ;
  		snc:cell_measures = "area: areacella" ;
  		snc:history = "2012-05-18T15:38:52Z altered by CMOR: replaced missing value flag (1e+36) with standard missing value (1e+20)." ;
  		snc:missing_value = 1.e+20f ;
  		snc:_FillValue = 1.e+20f ;
  		snc:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_landIce_fx_CESM1-CAM5_historical_r0i0p0.nc areacella: areacella_fx_CESM1-CAM5_historical_r0i0p0.nc" ;
  	double time(time) ;
  		time:bounds = "time_bnds" ;
  		time:units = "days since 1850-01-01 00:00:00" ;
  		time:calendar = "noleap" ;
  		time:axis = "T" ;
  		time:long_name = "time" ;
  		time:standard_name = "time" ;
  	double time_bnds(time, bnds) ;

  // group attributes:
  		:institution = "NSF/DOE NCAR (National Center for Atmospheric Research) Boulder, CO, USA" ;
  		:institute_id = "NSF-DOE-NCAR" ;
  		:experiment_id = "historical" ;
  		:source = "CESM1-CAM5" ;
  		:model_id = "CESM1-CAM5" ;
  		:forcing = "Sl GHG Vl SS Ds SD BC MD OC Oz AA LU" ;
  		:parent_experiment_id = "piControl" ;
  		:parent_experiment_rip = "r1i1p1" ;
  		:branch_time = 2. ;
  		:contact = "cesm_data@ucar.edu" ;
  		:comment = "CESM home page: http://www.cesm.ucar.edu" ;
  		:references = "Neale, R., et.al. 2012: Coupled simulations from CESM1 using the Community Atmosphere Model version 5: (CAM5). See also http://www.cesm.ucar.edu/publications" ;
  		:initialization_method = 1 ;
  		:physics_version = 1 ;
  		:tracking_id = "2ee6c8fd-9752-4455-bed3-576a01e9fed6" ;
  		:acknowledgements = "The CESM project is supported by the National Science Foundation and the Office of Science (BER) of the U.S. Department of Energy. NCAR is sponsored by the National Science Foundation. This research used resources of the Oak Ridge Leadership Computing Facility, located in the National Center for Computational Sciences at Oak Ridge National Laboratory, which is supported by the Office of Science (BER) of the Department of Energy under Contract DE-AC05-00OR22725." ;
  		:cesm_casename = "b40_20th_1d_b08c5cn_138j" ;
  		:cesm_repotag = "cesm1_0_beta08" ;
  		:cesm_compset = "B20TRC5CN" ;
  		:resolution = "f09_g16 (0.9x1.25_gx1v6)" ;
  		:forcing_note = "Additional information on the external forcings used in this experiment can be found at http://www.cesm.ucar.edu/CMIP5/forcing_information" ;
  		:processed_by = "strandwg on silver.cgd.ucar.edu at 20120518  -093852.130" ;
  		:processing_code_information = "Last Changed Rev: 776 Last Changed Date: 2012-05-17 09:36:52 -0600 (Thu, 17 May 2012) Repository UUID: d2181dbe-5796-6825-dc7f-cbd98591f93d" ;
  		:product = "output" ;
  		:experiment = "historical" ;
  		:frequency = "mon" ;
  		:creation_date = "2012-05-18T15:38:54Z" ;
  		:history = "Sun Dec 30 19:53:35 2012: ncks -d time,1990-01-01 00:00:0.0, /media/grele_data/wenshan/cesm/historical-exp/snc_LImon_CESM1-CAM5_historical_r1i1p1_185001-200512.nc /media/grele_data/wenshan/cesm/historical-exp/snc_LImon_CESM1-CAM5_historical_r1i1p1_199001-200512.nc\n2012-05-18T15:38:54Z CMOR rewrote data to comply with CF standards and CMIP5 requirements." ;
  		:Conventions = "CF-1.4" ;
  		:project_id = "CMIP5" ;
  		:table_id = "Table LImon (12 January 2012) 429410275cb5466e41180ad9466db1bf" ;
  		:title = "CESM1-CAM5 model output prepared for CMIP5 historical" ;
  		:parent_experiment = "pre-industrial control" ;
  		:modeling_realm = "landIce land" ;
  		:realization = 1 ;
  		:cmor_version = "2.8.1" ;
  		:NCO = "20121231" ;
  data:

   lat = 0 ;

   lat_bnds = -0.46875, 0.46875 ;

   lon = 179.375 ;

   lon_bnds = 178.752170138889, 180 ;

   snc = 62.07145, 60.97509, 57.9104, 53.65452, 46.13708, 39.71951, 34.45684, 
      33.34816, 36.30897, 45.20145, 54.7042, 60.06191, 61.81068, 61.57235, 
      58.69954, 53.0875, 44.43778, 38.41296, 33.89512, 33.16334, 35.38866, 
      44.20527, 55.24973, 60.42582, 61.78408, 60.30222, 57.74767, 51.87217, 
      45.43856, 39.859, 34.65273, 33.69739, 35.79815, 45.94585, 55.98174, 
      60.11427, 62.11591, 61.35354, 58.43501, 52.39944, 45.27255, 38.83994, 
      34.82337, 33.47124, 35.81379, 46.57481, 54.41116, 60.62625, 62.25172, 
      61.1827, 58.42628, 52.6358, 45.15274, 38.88607, 33.73675, 33.29869, 
      35.76462, 43.97408, 55.61646, 60.97946, 62.00888, 60.70457, 57.56046, 
      51.62181, 45.01118, 38.69769, 33.83691, 33.11338, 35.41447, 44.51177, 
      54.35133, 59.83762, 61.02993, 61.28046, 58.4234, 52.3585, 45.51928, 
      39.02513, 34.5911, 33.34881, 35.93228, 45.4144, 53.66666, 59.19072, 
      62.61044, 60.99728, 58.37831, 53.53175, 46.06737, 38.39714, 34.13896, 
      33.22199, 35.57574, 45.33149, 55.18364, 60.08348, 62.00661, 60.72526, 
      58.49016, 52.98635, 45.39072, 39.37619, 34.2319, 33.21686, 35.65197, 
      46.41065, 54.66462, 60.34342, 61.5855, 60.53594, 58.07879, 53.05131, 
      45.6369, 38.99934, 33.72679, 33.10427, 34.7771, 44.55233, 55.62511, 
      59.83138, 61.37432, 60.32346, 57.32902, 52.26272, 45.0841, 38.28241, 
      33.7456, 33.1823, 35.83283, 45.20584, 54.09948, 60.86015, 62.31863, 
      61.09036, 58.49607, 52.52017, 45.4707, 39.66387, 34.60744, 33.46476, 
      36.29692, 47.46539, 54.06594, 59.21001, 61.56113, 61.5031, 58.06651, 
      52.88129, 45.14191, 38.97267, 33.80598, 33.34988, 36.13751, 45.83525, 
      54.13206, 59.95444, 61.17745, 60.35199, 58.45913, 52.94626, 45.55574, 
      38.65861, 33.37043, 32.96347, 35.39613, 46.5092, 55.11117, 58.78823, 
      61.00055, 60.24277, 57.43545, 52.00771, 45.43082, 39.07673, 33.98228, 
      32.92905, 35.72621, 45.6367, 55.0639, 60.17884, 62.44907, 61.56859, 
      58.70348, 51.78551, 44.38303, 38.12561, 34.06507, 32.99229, 35.49913, 
      46.25829, 54.67482, 61.06555 ;

   time = 51115.5, 51145, 51174.5, 51205, 51235.5, 51266, 51296.5, 51327.5, 
      51358, 51388.5, 51419, 51449.5, 51480.5, 51510, 51539.5, 51570, 
      51600.5, 51631, 51661.5, 51692.5, 51723, 51753.5, 51784, 51814.5, 
      51845.5, 51875, 51904.5, 51935, 51965.5, 51996, 52026.5, 52057.5, 
      52088, 52118.5, 52149, 52179.5, 52210.5, 52240, 52269.5, 52300, 
      52330.5, 52361, 52391.5, 52422.5, 52453, 52483.5, 52514, 52544.5, 
      52575.5, 52605, 52634.5, 52665, 52695.5, 52726, 52756.5, 52787.5, 
      52818, 52848.5, 52879, 52909.5, 52940.5, 52970, 52999.5, 53030, 
      53060.5, 53091, 53121.5, 53152.5, 53183, 53213.5, 53244, 53274.5, 
      53305.5, 53335, 53364.5, 53395, 53425.5, 53456, 53486.5, 53517.5, 
      53548, 53578.5, 53609, 53639.5, 53670.5, 53700, 53729.5, 53760, 
      53790.5, 53821, 53851.5, 53882.5, 53913, 53943.5, 53974, 54004.5, 
      54035.5, 54065, 54094.5, 54125, 54155.5, 54186, 54216.5, 54247.5, 
      54278, 54308.5, 54339, 54369.5, 54400.5, 54430, 54459.5, 54490, 
      54520.5, 54551, 54581.5, 54612.5, 54643, 54673.5, 54704, 54734.5, 
      54765.5, 54795, 54824.5, 54855, 54885.5, 54916, 54946.5, 54977.5, 
      55008, 55038.5, 55069, 55099.5, 55130.5, 55160, 55189.5, 55220, 
      55250.5, 55281, 55311.5, 55342.5, 55373, 55403.5, 55434, 55464.5, 
      55495.5, 55525, 55554.5, 55585, 55615.5, 55646, 55676.5, 55707.5, 
      55738, 55768.5, 55799, 55829.5, 55860.5, 55890, 55919.5, 55950, 
      55980.5, 56011, 56041.5, 56072.5, 56103, 56133.5, 56164, 56194.5, 
      56225.5, 56255, 56284.5, 56315, 56345.5, 56376, 56406.5, 56437.5, 
      56468, 56498.5, 56529, 56559.5, 56590.5, 56620, 56649.5, 56680, 
      56710.5, 56741, 56771.5, 56802.5, 56833, 56863.5, 56894, 56924.5 ;

   time_bnds =
  51100, 51131,
  51131, 51159,
  51159, 51190,
  51190, 51220,
  51220, 51251,
  51251, 51281,
  51281, 51312,
  51312, 51343,
  51343, 51373,
  51373, 51404,
  51404, 51434,
  51434, 51465,
  51465, 51496,
  51496, 51524,
  51524, 51555,
  51555, 51585,
  51585, 51616,
  51616, 51646,
  51646, 51677,
  51677, 51708,
  51708, 51738,
  51738, 51769,
  51769, 51799,
  51799, 51830,
  51830, 51861,
  51861, 51889,
  51889, 51920,
  51920, 51950,
  51950, 51981,
  51981, 52011,
  52011, 52042,
  52042, 52073,
  52073, 52103,
  52103, 52134,
  52134, 52164,
  52164, 52195,
  52195, 52226,
  52226, 52254,
  52254, 52285,
  52285, 52315,
  52315, 52346,
  52346, 52376,
  52376, 52407,
  52407, 52438,
  52438, 52468,
  52468, 52499,
  52499, 52529,
  52529, 52560,
  52560, 52591,
  52591, 52619,
  52619, 52650,
  52650, 52680,
  52680, 52711,
  52711, 52741,
  52741, 52772,
  52772, 52803,
  52803, 52833,
  52833, 52864,
  52864, 52894,
  52894, 52925,
  52925, 52956,
  52956, 52984,
  52984, 53015,
  53015, 53045,
  53045, 53076,
  53076, 53106,
  53106, 53137,
  53137, 53168,
  53168, 53198,
  53198, 53229,
  53229, 53259,
  53259, 53290,
  53290, 53321,
  53321, 53349,
  53349, 53380,
  53380, 53410,
  53410, 53441,
  53441, 53471,
  53471, 53502,
  53502, 53533,
  53533, 53563,
  53563, 53594,
  53594, 53624,
  53624, 53655,
  53655, 53686,
  53686, 53714,
  53714, 53745,
  53745, 53775,
  53775, 53806,
  53806, 53836,
  53836, 53867,
  53867, 53898,
  53898, 53928,
  53928, 53959,
  53959, 53989,
  53989, 54020,
  54020, 54051,
  54051, 54079,
  54079, 54110,
  54110, 54140,
  54140, 54171,
  54171, 54201,
  54201, 54232,
  54232, 54263,
  54263, 54293,
  54293, 54324,
  54324, 54354,
  54354, 54385,
  54385, 54416,
  54416, 54444,
  54444, 54475,
  54475, 54505,
  54505, 54536,
  54536, 54566,
  54566, 54597,
  54597, 54628,
  54628, 54658,
  54658, 54689,
  54689, 54719,
  54719, 54750,
  54750, 54781,
  54781, 54809,
  54809, 54840,
  54840, 54870,
  54870, 54901,
  54901, 54931,
  54931, 54962,
  54962, 54993,
  54993, 55023,
  55023, 55054,
  55054, 55084,
  55084, 55115,
  55115, 55146,
  55146, 55174,
  55174, 55205,
  55205, 55235,
  55235, 55266,
  55266, 55296,
  55296, 55327,
  55327, 55358,
  55358, 55388,
  55388, 55419,
  55419, 55449,
  55449, 55480,
  55480, 55511,
  55511, 55539,
  55539, 55570,
  55570, 55600,
  55600, 55631,
  55631, 55661,
  55661, 55692,
  55692, 55723,
  55723, 55753,
  55753, 55784,
  55784, 55814,
  55814, 55845,
  55845, 55876,
  55876, 55904,
  55904, 55935,
  55935, 55965,
  55965, 55996,
  55996, 56026,
  56026, 56057,
  56057, 56088,
  56088, 56118,
  56118, 56149,
  56149, 56179,
  56179, 56210,
  56210, 56241,
  56241, 56269,
  56269, 56300,
  56300, 56330,
  56330, 56361,
  56361, 56391,
  56391, 56422,
  56422, 56453,
  56453, 56483,
  56483, 56514,
  56514, 56544,
  56544, 56575,
  56575, 56606,
  56606, 56634,
  56634, 56665,
  56665, 56695,
  56695, 56726,
  56726, 56756,
  56756, 56787,
  56787, 56818,
  56818, 56848,
  56848, 56879,
  56879, 56909,
  56909, 56940 ;
  } // group snc_LImon_CESM1-CAM5_historical_r1i1p1_199001-200512

group: snc_LImon_CESM1-FASTCHEM_historical_r1i1p1_199001-200512 {
  dimensions:
  	bnds = 2 ;
  	time = 192 ;
  variables:
  	double lat ;
  		lat:bounds = "lat_bnds" ;
  		lat:units = "degrees_north" ;
  		lat:axis = "Y" ;
  		lat:long_name = "latitude" ;
  		lat:standard_name = "latitude" ;
  	double lat_bnds(bnds) ;
  	double lon ;
  		lon:bounds = "lon_bnds" ;
  		lon:units = "degrees_east" ;
  		lon:axis = "X" ;
  		lon:long_name = "longitude" ;
  		lon:standard_name = "longitude" ;
  	double lon_bnds(bnds) ;
  	float snc(time) ;
  		snc:standard_name = "surface_snow_area_fraction" ;
  		snc:long_name = "Snow Area Fraction" ;
  		snc:comment = "FSNO, CMIP5_table_comment: Fraction of each grid cell that is occupied by snow that rests on land portion of cell." ;
  		snc:units = "%" ;
  		snc:original_name = "FSNO" ;
  		snc:cell_methods = "time: mean (interval: 30 days)" ;
  		snc:cell_measures = "area: areacella" ;
  		snc:history = "2012-05-17T14:29:14Z altered by CMOR: replaced missing value flag (1e+36) with standard missing value (1e+20)." ;
  		snc:missing_value = 1.e+20f ;
  		snc:_FillValue = 1.e+20f ;
  		snc:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_landIce_fx_CESM1-FASTCHEM_historical_r0i0p0.nc areacella: areacella_fx_CESM1-FASTCHEM_historical_r0i0p0.nc" ;
  	double time(time) ;
  		time:bounds = "time_bnds" ;
  		time:units = "days since 1850-01-01 00:00:00" ;
  		time:calendar = "noleap" ;
  		time:axis = "T" ;
  		time:long_name = "time" ;
  		time:standard_name = "time" ;
  	double time_bnds(time, bnds) ;

  // group attributes:
  		:institution = "NSF/DOE NCAR (National Center for Atmospheric Research) Boulder, CO, USA" ;
  		:institute_id = "NSF-DOE-NCAR" ;
  		:experiment_id = "historical" ;
  		:source = "CESM1-FASTCHEM" ;
  		:model_id = "CESM1-FASTCHEM" ;
  		:forcing = "Sl GHG Vl SS Ds SD BC MD OC Oz AA LU" ;
  		:parent_experiment_id = "piControl" ;
  		:parent_experiment_rip = "r1i1p1" ;
  		:branch_time = 0. ;
  		:contact = "cesm_data@ucar.edu" ;
  		:comment = "CESM home page: http://www.cesm.ucar.edu" ;
  		:references = "TBD" ;
  		:initialization_method = 1 ;
  		:physics_version = 1 ;
  		:tracking_id = "6b2ee7c3-9fd1-41e8-81d3-363f5f40b846" ;
  		:acknowledgements = "The CESM project is supported by the National Science Foundation and the Office of Science (BER) of the U.S. Department of Energy. NCAR is sponsored by the National Science Foundation. Computing resources were provided by the Climate Simulation Laboratory at the NCAR Computational and Information Systems Laboratory (CISL), sponsored by the National Science Foundation and other agencies." ;
  		:cesm_casename = "b40.20th.1deg.fschem.002" ;
  		:cesm_repotag = "ccsm4_0_beta55" ;
  		:cesm_compset = "B20TRCNCHM" ;
  		:resolution = "f09_g16 (0.9x1.25_gx1v6)" ;
  		:forcing_note = "Additional information on the external forcings used in this experiment can be found at http://www.cesm.ucar.edu/CMIP5/forcing_information" ;
  		:processed_by = "strandwg on silver.cgd.ucar.edu at 20120517  -082914.590" ;
  		:processing_code_information = "Last Changed Rev: 774 Last Changed Date: 2012-05-16 16:39:53 -0600 (Wed, 16 May 2012) Repository UUID: d2181dbe-5796-6825-dc7f-cbd98591f93d" ;
  		:product = "output" ;
  		:experiment = "historical" ;
  		:frequency = "mon" ;
  		:creation_date = "2012-05-17T14:29:16Z" ;
  		:history = "Sun Dec 30 18:44:33 2012: ncks -d time,1990-01-01 00:00:0.0, /media/grele_data/wenshan/cesm/atmos-his/snc_LImon_CESM1-FASTCHEM_historical_r1i1p1_185001-200512.nc /media/grele_data/wenshan/cesm/atmos-his/snc_LImon_CESM1-FASTCHEM_historical_r1i1p1_199001-200512.nc\n2012-05-17T14:29:16Z CMOR rewrote data to comply with CF standards and CMIP5 requirements." ;
  		:Conventions = "CF-1.4" ;
  		:project_id = "CMIP5" ;
  		:table_id = "Table LImon (12 January 2012) 429410275cb5466e41180ad9466db1bf" ;
  		:title = "CESM1-FASTCHEM model output prepared for CMIP5 historical" ;
  		:parent_experiment = "pre-industrial control" ;
  		:modeling_realm = "landIce land" ;
  		:realization = 1 ;
  		:cmor_version = "2.8.1" ;
  		:NCO = "20121231" ;
  data:

   lat = 0 ;

   lat_bnds = -0.46875, 0.46875 ;

   lon = 179.375 ;

   lon_bnds = 178.752170138889, 180 ;

   snc = 61.35922, 60.11757, 56.77606, 51.86809, 44.5789, 38.14515, 33.07576, 
      33.10382, 36.08701, 44.22195, 53.31831, 58.38189, 61.49045, 61.94424, 
      57.49084, 51.4422, 45.94965, 39.01295, 33.63499, 32.85659, 37.11253, 
      44.66447, 53.68621, 59.86607, 60.47795, 60.76228, 56.93726, 51.28774, 
      44.71006, 38.61081, 33.86168, 33.20221, 36.73127, 47.33617, 56.14992, 
      59.57047, 61.68317, 60.56863, 57.71325, 52.03714, 45.42717, 37.95629, 
      34.18681, 33.22436, 37.29691, 46.26162, 54.90151, 60.79268, 61.64498, 
      61.18701, 58.2198, 51.28855, 44.98966, 38.63614, 33.35585, 32.91083, 
      36.14466, 44.34061, 55.25936, 59.61454, 60.81066, 59.89703, 56.78886, 
      51.34318, 44.89197, 37.97543, 33.65519, 32.92331, 34.96158, 46.80618, 
      54.58622, 60.04884, 62.42439, 61.58648, 58.25958, 52.32566, 44.83265, 
      37.18033, 33.52879, 33.03136, 36.15388, 46.12405, 53.96253, 59.95536, 
      60.54895, 58.84748, 56.34169, 50.48568, 43.52483, 38.12297, 33.95269, 
      33.15511, 35.92193, 43.6329, 54.4885, 58.7534, 59.50955, 59.38222, 
      56.4384, 50.68229, 44.19793, 37.82106, 33.37074, 33.17641, 36.68989, 
      44.85901, 53.11116, 57.75417, 60.42802, 59.57334, 56.00442, 50.08305, 
      43.97726, 38.49365, 33.53299, 32.87168, 35.67901, 45.14764, 53.06521, 
      58.36853, 60.57628, 59.72157, 56.75367, 50.25916, 43.97816, 38.27824, 
      33.78714, 33.07768, 35.71507, 43.82384, 53.86621, 59.8281, 62.98288, 
      60.35318, 56.95187, 50.56234, 44.47134, 37.65242, 33.04737, 32.78938, 
      35.73754, 45.56456, 53.15977, 58.71597, 59.50213, 59.8814, 57.11369, 
      51.297, 45.74558, 38.31946, 33.30605, 32.88755, 35.60548, 43.45373, 
      53.75446, 58.68278, 59.57464, 59.02721, 56.63763, 51.11911, 43.58306, 
      36.49274, 33.1369, 32.70171, 35.42366, 45.84877, 52.81328, 58.69426, 
      60.35154, 58.81255, 56.24924, 51.00918, 44.1529, 38.16121, 33.06249, 
      32.81034, 35.65083, 44.37822, 52.15639, 59.87329, 61.16865, 60.83504, 
      56.66895, 51.41212, 43.97941, 37.59834, 33.35089, 32.66173, 34.87273, 
      44.44268, 52.47154, 58.85749 ;

   time = 51115.5, 51145, 51174.5, 51205, 51235.5, 51266, 51296.5, 51327.5, 
      51358, 51388.5, 51419, 51449.5, 51480.5, 51510, 51539.5, 51570, 
      51600.5, 51631, 51661.5, 51692.5, 51723, 51753.5, 51784, 51814.5, 
      51845.5, 51875, 51904.5, 51935, 51965.5, 51996, 52026.5, 52057.5, 
      52088, 52118.5, 52149, 52179.5, 52210.5, 52240, 52269.5, 52300, 
      52330.5, 52361, 52391.5, 52422.5, 52453, 52483.5, 52514, 52544.5, 
      52575.5, 52605, 52634.5, 52665, 52695.5, 52726, 52756.5, 52787.5, 
      52818, 52848.5, 52879, 52909.5, 52940.5, 52970, 52999.5, 53030, 
      53060.5, 53091, 53121.5, 53152.5, 53183, 53213.5, 53244, 53274.5, 
      53305.5, 53335, 53364.5, 53395, 53425.5, 53456, 53486.5, 53517.5, 
      53548, 53578.5, 53609, 53639.5, 53670.5, 53700, 53729.5, 53760, 
      53790.5, 53821, 53851.5, 53882.5, 53913, 53943.5, 53974, 54004.5, 
      54035.5, 54065, 54094.5, 54125, 54155.5, 54186, 54216.5, 54247.5, 
      54278, 54308.5, 54339, 54369.5, 54400.5, 54430, 54459.5, 54490, 
      54520.5, 54551, 54581.5, 54612.5, 54643, 54673.5, 54704, 54734.5, 
      54765.5, 54795, 54824.5, 54855, 54885.5, 54916, 54946.5, 54977.5, 
      55008, 55038.5, 55069, 55099.5, 55130.5, 55160, 55189.5, 55220, 
      55250.5, 55281, 55311.5, 55342.5, 55373, 55403.5, 55434, 55464.5, 
      55495.5, 55525, 55554.5, 55585, 55615.5, 55646, 55676.5, 55707.5, 
      55738, 55768.5, 55799, 55829.5, 55860.5, 55890, 55919.5, 55950, 
      55980.5, 56011, 56041.5, 56072.5, 56103, 56133.5, 56164, 56194.5, 
      56225.5, 56255, 56284.5, 56315, 56345.5, 56376, 56406.5, 56437.5, 
      56468, 56498.5, 56529, 56559.5, 56590.5, 56620, 56649.5, 56680, 
      56710.5, 56741, 56771.5, 56802.5, 56833, 56863.5, 56894, 56924.5 ;

   time_bnds =
  51100, 51131,
  51131, 51159,
  51159, 51190,
  51190, 51220,
  51220, 51251,
  51251, 51281,
  51281, 51312,
  51312, 51343,
  51343, 51373,
  51373, 51404,
  51404, 51434,
  51434, 51465,
  51465, 51496,
  51496, 51524,
  51524, 51555,
  51555, 51585,
  51585, 51616,
  51616, 51646,
  51646, 51677,
  51677, 51708,
  51708, 51738,
  51738, 51769,
  51769, 51799,
  51799, 51830,
  51830, 51861,
  51861, 51889,
  51889, 51920,
  51920, 51950,
  51950, 51981,
  51981, 52011,
  52011, 52042,
  52042, 52073,
  52073, 52103,
  52103, 52134,
  52134, 52164,
  52164, 52195,
  52195, 52226,
  52226, 52254,
  52254, 52285,
  52285, 52315,
  52315, 52346,
  52346, 52376,
  52376, 52407,
  52407, 52438,
  52438, 52468,
  52468, 52499,
  52499, 52529,
  52529, 52560,
  52560, 52591,
  52591, 52619,
  52619, 52650,
  52650, 52680,
  52680, 52711,
  52711, 52741,
  52741, 52772,
  52772, 52803,
  52803, 52833,
  52833, 52864,
  52864, 52894,
  52894, 52925,
  52925, 52956,
  52956, 52984,
  52984, 53015,
  53015, 53045,
  53045, 53076,
  53076, 53106,
  53106, 53137,
  53137, 53168,
  53168, 53198,
  53198, 53229,
  53229, 53259,
  53259, 53290,
  53290, 53321,
  53321, 53349,
  53349, 53380,
  53380, 53410,
  53410, 53441,
  53441, 53471,
  53471, 53502,
  53502, 53533,
  53533, 53563,
  53563, 53594,
  53594, 53624,
  53624, 53655,
  53655, 53686,
  53686, 53714,
  53714, 53745,
  53745, 53775,
  53775, 53806,
  53806, 53836,
  53836, 53867,
  53867, 53898,
  53898, 53928,
  53928, 53959,
  53959, 53989,
  53989, 54020,
  54020, 54051,
  54051, 54079,
  54079, 54110,
  54110, 54140,
  54140, 54171,
  54171, 54201,
  54201, 54232,
  54232, 54263,
  54263, 54293,
  54293, 54324,
  54324, 54354,
  54354, 54385,
  54385, 54416,
  54416, 54444,
  54444, 54475,
  54475, 54505,
  54505, 54536,
  54536, 54566,
  54566, 54597,
  54597, 54628,
  54628, 54658,
  54658, 54689,
  54689, 54719,
  54719, 54750,
  54750, 54781,
  54781, 54809,
  54809, 54840,
  54840, 54870,
  54870, 54901,
  54901, 54931,
  54931, 54962,
  54962, 54993,
  54993, 55023,
  55023, 55054,
  55054, 55084,
  55084, 55115,
  55115, 55146,
  55146, 55174,
  55174, 55205,
  55205, 55235,
  55235, 55266,
  55266, 55296,
  55296, 55327,
  55327, 55358,
  55358, 55388,
  55388, 55419,
  55419, 55449,
  55449, 55480,
  55480, 55511,
  55511, 55539,
  55539, 55570,
  55570, 55600,
  55600, 55631,
  55631, 55661,
  55661, 55692,
  55692, 55723,
  55723, 55753,
  55753, 55784,
  55784, 55814,
  55814, 55845,
  55845, 55876,
  55876, 55904,
  55904, 55935,
  55935, 55965,
  55965, 55996,
  55996, 56026,
  56026, 56057,
  56057, 56088,
  56088, 56118,
  56118, 56149,
  56149, 56179,
  56179, 56210,
  56210, 56241,
  56241, 56269,
  56269, 56300,
  56300, 56330,
  56330, 56361,
  56361, 56391,
  56391, 56422,
  56422, 56453,
  56453, 56483,
  56483, 56514,
  56514, 56544,
  56544, 56575,
  56575, 56606,
  56606, 56634,
  56634, 56665,
  56665, 56695,
  56695, 56726,
  56726, 56756,
  56756, 56787,
  56787, 56818,
  56818, 56848,
  56848, 56879,
  56879, 56909,
  56909, 56940 ;
  } // group snc_LImon_CESM1-FASTCHEM_historical_r1i1p1_199001-200512

group: snc_LImon_CESM1-WACCM_historical_r1i1p1_199001-200512 {
  dimensions:
  	bnds = 2 ;
  	time = 192 ;
  variables:
  	double lat ;
  		lat:bounds = "lat_bnds" ;
  		lat:units = "degrees_north" ;
  		lat:axis = "Y" ;
  		lat:long_name = "latitude" ;
  		lat:standard_name = "latitude" ;
  	double lat_bnds(bnds) ;
  	double lon ;
  		lon:bounds = "lon_bnds" ;
  		lon:units = "degrees_east" ;
  		lon:axis = "X" ;
  		lon:long_name = "longitude" ;
  		lon:standard_name = "longitude" ;
  	double lon_bnds(bnds) ;
  	float snc(time) ;
  		snc:standard_name = "surface_snow_area_fraction" ;
  		snc:long_name = "Snow Area Fraction" ;
  		snc:comment = "FSNO, CMIP5_table_comment: Fraction of each grid cell that is occupied by snow that rests on land portion of cell." ;
  		snc:units = "%" ;
  		snc:original_name = "FSNO" ;
  		snc:cell_methods = "time: mean (interval: 30 days)" ;
  		snc:cell_measures = "area: areacella" ;
  		snc:history = "2012-05-31T13:28:20Z altered by CMOR: replaced missing value flag (1e+36) with standard missing value (1e+20)." ;
  		snc:missing_value = 1.e+20f ;
  		snc:_FillValue = 1.e+20f ;
  		snc:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_landIce_fx_CESM1-WACCM_historical_r0i0p0.nc areacella: areacella_fx_CESM1-WACCM_historical_r0i0p0.nc" ;
  	double time(time) ;
  		time:bounds = "time_bnds" ;
  		time:units = "days since 1850-01-01 00:00:00" ;
  		time:calendar = "noleap" ;
  		time:axis = "T" ;
  		time:long_name = "time" ;
  		time:standard_name = "time" ;
  	double time_bnds(time, bnds) ;

  // group attributes:
  		:institution = "NSF/DOE NCAR (National Center for Atmospheric Research) Boulder, CO, USA" ;
  		:institute_id = "NSF-DOE-NCAR" ;
  		:experiment_id = "historical" ;
  		:source = "CESM1-WACCM" ;
  		:model_id = "CESM1-WACCM" ;
  		:forcing = "Sl GHG Vl SS Ds SD BC MD OC Oz AA LU" ;
  		:parent_experiment_id = "piControl" ;
  		:parent_experiment_rip = "r1i1p1" ;
  		:branch_time = 1. ;
  		:contact = "cesm_data@ucar.edu" ;
  		:comment = "CESM home page: http://www.cesm.ucar.edu" ;
  		:references = "Marsh, D., et.al. 2012: WACCM4 simulations of atmospheric trends from 1850 to present. See also http://www.cesm.ucar.edu/publications" ;
  		:initialization_method = 1 ;
  		:physics_version = 1 ;
  		:tracking_id = "ef93cac6-c5d8-4b32-9ff0-9cbd27d8e66a" ;
  		:acknowledgements = "The CESM project is supported by the National Science Foundation and the Office of Science (BER) of the U.S. Department of Energy. NCAR is sponsored by the National Science Foundation. Computing resources were provided by the Climate Simulation Laboratory at the NCAR Computational and Information Systems Laboratory (CISL), sponsored by the National Science Foundation and other agencies." ;
  		:cesm_casename = "b40.20th.track1.2deg.wcm.007" ;
  		:cesm_repotag = "ccsm4_0_beta52" ;
  		:cesm_compset = "BW20TRCN" ;
  		:resolution = "f19_g16 (1.9x2.5_gx1v6)" ;
  		:forcing_note = "Additional information on the external forcings used in this experiment can be found at http://www.cesm.ucar.edu/CMIP5/forcing_information" ;
  		:processed_by = "strandwg on mirage3 at 20120531  -072820.637" ;
  		:processing_code_information = "Last Changed Rev: 820 Last Changed Date: 2012-05-30 15:07:51 -0600 (Wed, 30 May 2012) Repository UUID: d2181dbe-5796-6825-dc7f-cbd98591f93d" ;
  		:product = "output" ;
  		:experiment = "historical" ;
  		:frequency = "mon" ;
  		:creation_date = "2012-05-31T13:28:21Z" ;
  		:history = "Sun Dec 30 18:44:48 2012: ncks -d time,1990-01-01 00:00:0.0, /media/grele_data/wenshan/cesm/atmos-his/snc_LImon_CESM1-WACCM_historical_r1i1p1_185001-200512.nc /media/grele_data/wenshan/cesm/atmos-his/snc_LImon_CESM1-WACCM_historical_r1i1p1_199001-200512.nc\n2012-05-31T13:28:21Z CMOR rewrote data to comply with CF standards and CMIP5 requirements." ;
  		:Conventions = "CF-1.4" ;
  		:project_id = "CMIP5" ;
  		:table_id = "Table LImon (12 January 2012) 429410275cb5466e41180ad9466db1bf" ;
  		:title = "CESM1-WACCM model output prepared for CMIP5 historical" ;
  		:parent_experiment = "pre-industrial control" ;
  		:modeling_realm = "landIce land" ;
  		:realization = 1 ;
  		:cmor_version = "2.8.1" ;
  		:NCO = "20121231" ;
  data:

   lat = 0 ;

   lat_bnds = -0.9375, 0.9375 ;

   lon = 178.75 ;

   lon_bnds = 177.508680555556, 180 ;

   snc = 58.30264, 57.57164, 55.40315, 51.30324, 44.92303, 38.5704, 34.73244, 
      33.40054, 36.39927, 44.70775, 52.15816, 56.68031, 58.03102, 57.54689, 
      55.26139, 50.4637, 43.77814, 37.38792, 33.62425, 33.55622, 36.64553, 
      45.27554, 52.15833, 58.00319, 60.39744, 60.92056, 57.63554, 49.88797, 
      43.92668, 38.43521, 34.53812, 33.3124, 35.9039, 44.06456, 52.36027, 
      57.0512, 58.79975, 58.51964, 56.20938, 51.16467, 44.37978, 36.94592, 
      33.22895, 33.14706, 36.17453, 45.27049, 52.18351, 57.12118, 59.51681, 
      58.67272, 55.35041, 49.88683, 44.25735, 38.44041, 33.5755, 32.74223, 
      35.94821, 45.38294, 52.94146, 57.9625, 59.15063, 58.10602, 55.73347, 
      50.96825, 44.56723, 38.10284, 33.3599, 32.98213, 35.90267, 43.69198, 
      53.58926, 58.14558, 59.82616, 58.78763, 56.74655, 51.95066, 45.35992, 
      36.72455, 32.72494, 32.69721, 35.77222, 44.46194, 52.06679, 56.87531, 
      59.6659, 58.29536, 54.9007, 49.42334, 43.95756, 36.97405, 33.28221, 
      32.84733, 35.55394, 44.29796, 52.48971, 57.30995, 58.13997, 57.98017, 
      55.87465, 50.05117, 43.26404, 36.44524, 33.10003, 32.76156, 35.33764, 
      43.94565, 51.96738, 57.09196, 58.89738, 58.25306, 56.59516, 52.6945, 
      44.78914, 37.78814, 32.69427, 32.55199, 36.63308, 45.10502, 52.95998, 
      58.76827, 60.31608, 58.63898, 56.55276, 51.78586, 44.54252, 37.68716, 
      33.18846, 32.67733, 35.96641, 44.42927, 52.38469, 57.34024, 58.62802, 
      58.19473, 54.8047, 48.94669, 42.90043, 37.16561, 33.53363, 32.7061, 
      35.18901, 43.03574, 51.86749, 57.74329, 60.09589, 60.36689, 57.27032, 
      50.42865, 44.00283, 37.74604, 33.42166, 32.72996, 35.66089, 43.93026, 
      51.86792, 56.20585, 59.0007, 56.74605, 55.26267, 50.96566, 44.89715, 
      39.17544, 33.97953, 33.06948, 35.02919, 41.76595, 51.58342, 57.55459, 
      59.76404, 59.17727, 56.35314, 51.4416, 44.05042, 37.53273, 33.42004, 
      33.01108, 35.84677, 44.90015, 52.5538, 57.30947, 60.00209, 59.43186, 
      55.75416, 50.16666, 42.99211, 37.32963, 33.30409, 32.98776, 34.92936, 
      42.45069, 51.19328, 58.13653 ;

   time = 51115.5, 51145, 51174.5, 51205, 51235.5, 51266, 51296.5, 51327.5, 
      51358, 51388.5, 51419, 51449.5, 51480.5, 51510, 51539.5, 51570, 
      51600.5, 51631, 51661.5, 51692.5, 51723, 51753.5, 51784, 51814.5, 
      51845.5, 51875, 51904.5, 51935, 51965.5, 51996, 52026.5, 52057.5, 
      52088, 52118.5, 52149, 52179.5, 52210.5, 52240, 52269.5, 52300, 
      52330.5, 52361, 52391.5, 52422.5, 52453, 52483.5, 52514, 52544.5, 
      52575.5, 52605, 52634.5, 52665, 52695.5, 52726, 52756.5, 52787.5, 
      52818, 52848.5, 52879, 52909.5, 52940.5, 52970, 52999.5, 53030, 
      53060.5, 53091, 53121.5, 53152.5, 53183, 53213.5, 53244, 53274.5, 
      53305.5, 53335, 53364.5, 53395, 53425.5, 53456, 53486.5, 53517.5, 
      53548, 53578.5, 53609, 53639.5, 53670.5, 53700, 53729.5, 53760, 
      53790.5, 53821, 53851.5, 53882.5, 53913, 53943.5, 53974, 54004.5, 
      54035.5, 54065, 54094.5, 54125, 54155.5, 54186, 54216.5, 54247.5, 
      54278, 54308.5, 54339, 54369.5, 54400.5, 54430, 54459.5, 54490, 
      54520.5, 54551, 54581.5, 54612.5, 54643, 54673.5, 54704, 54734.5, 
      54765.5, 54795, 54824.5, 54855, 54885.5, 54916, 54946.5, 54977.5, 
      55008, 55038.5, 55069, 55099.5, 55130.5, 55160, 55189.5, 55220, 
      55250.5, 55281, 55311.5, 55342.5, 55373, 55403.5, 55434, 55464.5, 
      55495.5, 55525, 55554.5, 55585, 55615.5, 55646, 55676.5, 55707.5, 
      55738, 55768.5, 55799, 55829.5, 55860.5, 55890, 55919.5, 55950, 
      55980.5, 56011, 56041.5, 56072.5, 56103, 56133.5, 56164, 56194.5, 
      56225.5, 56255, 56284.5, 56315, 56345.5, 56376, 56406.5, 56437.5, 
      56468, 56498.5, 56529, 56559.5, 56590.5, 56620, 56649.5, 56680, 
      56710.5, 56741, 56771.5, 56802.5, 56833, 56863.5, 56894, 56924.5 ;

   time_bnds =
  51100, 51131,
  51131, 51159,
  51159, 51190,
  51190, 51220,
  51220, 51251,
  51251, 51281,
  51281, 51312,
  51312, 51343,
  51343, 51373,
  51373, 51404,
  51404, 51434,
  51434, 51465,
  51465, 51496,
  51496, 51524,
  51524, 51555,
  51555, 51585,
  51585, 51616,
  51616, 51646,
  51646, 51677,
  51677, 51708,
  51708, 51738,
  51738, 51769,
  51769, 51799,
  51799, 51830,
  51830, 51861,
  51861, 51889,
  51889, 51920,
  51920, 51950,
  51950, 51981,
  51981, 52011,
  52011, 52042,
  52042, 52073,
  52073, 52103,
  52103, 52134,
  52134, 52164,
  52164, 52195,
  52195, 52226,
  52226, 52254,
  52254, 52285,
  52285, 52315,
  52315, 52346,
  52346, 52376,
  52376, 52407,
  52407, 52438,
  52438, 52468,
  52468, 52499,
  52499, 52529,
  52529, 52560,
  52560, 52591,
  52591, 52619,
  52619, 52650,
  52650, 52680,
  52680, 52711,
  52711, 52741,
  52741, 52772,
  52772, 52803,
  52803, 52833,
  52833, 52864,
  52864, 52894,
  52894, 52925,
  52925, 52956,
  52956, 52984,
  52984, 53015,
  53015, 53045,
  53045, 53076,
  53076, 53106,
  53106, 53137,
  53137, 53168,
  53168, 53198,
  53198, 53229,
  53229, 53259,
  53259, 53290,
  53290, 53321,
  53321, 53349,
  53349, 53380,
  53380, 53410,
  53410, 53441,
  53441, 53471,
  53471, 53502,
  53502, 53533,
  53533, 53563,
  53563, 53594,
  53594, 53624,
  53624, 53655,
  53655, 53686,
  53686, 53714,
  53714, 53745,
  53745, 53775,
  53775, 53806,
  53806, 53836,
  53836, 53867,
  53867, 53898,
  53898, 53928,
  53928, 53959,
  53959, 53989,
  53989, 54020,
  54020, 54051,
  54051, 54079,
  54079, 54110,
  54110, 54140,
  54140, 54171,
  54171, 54201,
  54201, 54232,
  54232, 54263,
  54263, 54293,
  54293, 54324,
  54324, 54354,
  54354, 54385,
  54385, 54416,
  54416, 54444,
  54444, 54475,
  54475, 54505,
  54505, 54536,
  54536, 54566,
  54566, 54597,
  54597, 54628,
  54628, 54658,
  54658, 54689,
  54689, 54719,
  54719, 54750,
  54750, 54781,
  54781, 54809,
  54809, 54840,
  54840, 54870,
  54870, 54901,
  54901, 54931,
  54931, 54962,
  54962, 54993,
  54993, 55023,
  55023, 55054,
  55054, 55084,
  55084, 55115,
  55115, 55146,
  55146, 55174,
  55174, 55205,
  55205, 55235,
  55235, 55266,
  55266, 55296,
  55296, 55327,
  55327, 55358,
  55358, 55388,
  55388, 55419,
  55419, 55449,
  55449, 55480,
  55480, 55511,
  55511, 55539,
  55539, 55570,
  55570, 55600,
  55600, 55631,
  55631, 55661,
  55661, 55692,
  55692, 55723,
  55723, 55753,
  55753, 55784,
  55784, 55814,
  55814, 55845,
  55845, 55876,
  55876, 55904,
  55904, 55935,
  55935, 55965,
  55965, 55996,
  55996, 56026,
  56026, 56057,
  56057, 56088,
  56088, 56118,
  56118, 56149,
  56149, 56179,
  56179, 56210,
  56210, 56241,
  56241, 56269,
  56269, 56300,
  56300, 56330,
  56330, 56361,
  56361, 56391,
  56391, 56422,
  56422, 56453,
  56453, 56483,
  56483, 56514,
  56514, 56544,
  56544, 56575,
  56575, 56606,
  56606, 56634,
  56634, 56665,
  56665, 56695,
  56695, 56726,
  56726, 56756,
  56756, 56787,
  56787, 56818,
  56818, 56848,
  56848, 56879,
  56879, 56909,
  56909, 56940 ;
  } // group snc_LImon_CESM1-WACCM_historical_r1i1p1_199001-200512
}
