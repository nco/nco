// Generate netCDF file with:
// ncgen -k netCDF-4 -b -o ~/nco/data/obs.nc ~/nco/data/obs.cdl

netcdf obs {
  dimensions:
  time=4;
  variables:
  float tas(time);
  data:
  tas=273,273,273,273;
 
} // end root group
