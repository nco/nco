// $Header: /data/zender/nco_20150216/nco/bm/ipcc_dly_T85.cdl,v 1.1 2005-03-23 18:13:47 mangalam Exp $
// ncgen -b -o ipcc_dly_T85.nc ipcc_dly_T85.cdl (-> 1,142,957,636 bytes)
// takes about 48 (real) sec on 900MHz/512MB a22p thinkpad, 
// most of it waiting for disk

// Valid CDF/netCDF files need not have any defined variable or data
// Use ncap LHS-casting to define variables with big dimensions
netcdf ipcc_dly_T85{
dimensions:
    time=8;  // 'real' variables
    lev=32;
    lat=128;
    lon=256;
variables:
    double time(time);  // indices all have to be ints.
    double lev(lev);
    double lat(lat);
    double lon(lon);
    
// real variables
// 32 4D vars
    float d4_00(time,lev,lat,lon);
    float d4_01(time,lev,lat,lon);
    float d4_02(time,lev,lat,lon);
    float d4_03(time,lev,lat,lon);
    float d4_04(time,lev,lat,lon);
    float d4_05(time,lev,lat,lon);
    float d4_06(time,lev,lat,lon);
    float d4_07(time,lev,lat,lon);
    float d4_08(time,lev,lat,lon);
    float d4_09(time,lev,lat,lon);
    float d4_10(time,lev,lat,lon);
    float d4_11(time,lev,lat,lon);
    float d4_12(time,lev,lat,lon);
    float d4_13(time,lev,lat,lon);
    float d4_14(time,lev,lat,lon);
    float d4_15(time,lev,lat,lon);
    float d4_16(time,lev,lat,lon);
    float d4_17(time,lev,lat,lon);
    float d4_18(time,lev,lat,lon);
    float d4_19(time,lev,lat,lon);
    float d4_20(time,lev,lat,lon);
    float d4_21(time,lev,lat,lon);
    float d4_22(time,lev,lat,lon);
    float d4_23(time,lev,lat,lon);
    float d4_24(time,lev,lat,lon);
    float d4_25(time,lev,lat,lon);
    float d4_26(time,lev,lat,lon);
    float d4_27(time,lev,lat,lon);
    float d4_28(time,lev,lat,lon);
    float d4_29(time,lev,lat,lon);
    float d4_30(time,lev,lat,lon);
    float d4_31(time,lev,lat,lon);

//  64 3D vars
    float d3_00(time,lat,lon);
    float d3_01(time,lat,lon);
    float d3_02(time,lat,lon);
    float d3_03(time,lat,lon);
    float d3_04(time,lat,lon);
    float d3_05(time,lat,lon);
    float d3_06(time,lat,lon);
    float d3_07(time,lat,lon);
    float d3_08(time,lat,lon);
    float d3_09(time,lat,lon);
    float d3_10(time,lat,lon);
    float d3_11(time,lat,lon);
    float d3_12(time,lat,lon);
    float d3_13(time,lat,lon);
    float d3_14(time,lat,lon);
    float d3_15(time,lat,lon);
    float d3_16(time,lat,lon);
    float d3_17(time,lat,lon);
    float d3_18(time,lat,lon);
    float d3_19(time,lat,lon);
    float d3_20(time,lat,lon);
    float d3_21(time,lat,lon);
    float d3_22(time,lat,lon);
    float d3_23(time,lat,lon);
    float d3_24(time,lat,lon);
    float d3_25(time,lat,lon);
    float d3_26(time,lat,lon);
    float d3_27(time,lat,lon);
    float d3_28(time,lat,lon);
    float d3_29(time,lat,lon);
    float d3_30(time,lat,lon);
    float d3_31(time,lat,lon);
    float d3_32(time,lat,lon);
    float d3_33(time,lat,lon);
    float d3_34(time,lat,lon);
    float d3_35(time,lat,lon);
    float d3_36(time,lat,lon);
    float d3_37(time,lat,lon);
    float d3_38(time,lat,lon);
    float d3_39(time,lat,lon);
    float d3_40(time,lat,lon);
    float d3_41(time,lat,lon);
    float d3_42(time,lat,lon);
    float d3_43(time,lat,lon);
    float d3_44(time,lat,lon);
    float d3_45(time,lat,lon);
    float d3_46(time,lat,lon);
    float d3_47(time,lat,lon);
    float d3_48(time,lat,lon);
    float d3_49(time,lat,lon);
    float d3_50(time,lat,lon);
    float d3_51(time,lat,lon);
    float d3_52(time,lat,lon);
    float d3_53(time,lat,lon);
    float d3_54(time,lat,lon);
    float d3_55(time,lat,lon);
    float d3_56(time,lat,lon);
    float d3_57(time,lat,lon);
    float d3_58(time,lat,lon);
    float d3_59(time,lat,lon);
    float d3_60(time,lat,lon);
    float d3_61(time,lat,lon);
    float d3_62(time,lat,lon);
    float d3_63(time,lat,lon);

// 16 2D vars
    float d2_00(lat,lon);
    float d2_01(lat,lon);
    float d2_02(lat,lon);
    float d2_03(lat,lon);
    float d2_04(lat,lon);
    float d2_05(lat,lon);
    float d2_06(lat,lon);
    float d2_07(lat,lon);
    float d2_08(lat,lon);
    float d2_09(lat,lon);
    float d2_10(lat,lon);
    float d2_11(lat,lon);
    float d2_12(lat,lon);
    float d2_13(lat,lon);
    float d2_14(lat,lon);
    float d2_15(lat,lon);
    
// 8 1D vars
    float d1_00(time);
    float d1_01(time);
    float d1_02(time);
    float d1_03(time);
    float d1_04(time);
    float d1_05(time);
    float d1_06(time);
    float d1_07(time);

// 8 0D vars    
    float weepy;
    float dopey;
    float sleepy;
    float grouchy;
    float sneezy;
    float doc;
    float wanky;
    float skanky;

data:
    lat=0.703125,1.40625,2.109375,2.8125,3.515625,4.21875,4.921875,5.625,6.328125,7.03125,7.734375,8.4375,9.140625,9.84375,10.546875,11.25,11.953125,12.65625,13.359375,14.0625,14.765625,15.46875,16.171875,16.875,17.578125,18.28125,18.984375,19.6875,20.390625,21.09375,21.796875,22.5,23.203125,23.90625,24.609375,25.3125,26.015625,26.71875,27.421875,28.125,28.828125,29.53125,30.234375,30.9375,31.640625,32.34375,33.046875,33.75,34.453125,35.15625,35.859375,36.5625,37.265625,37.96875,38.671875,39.375,40.078125,40.78125,41.484375,42.1875,42.890625,43.59375,44.296875,45,45.703125,46.40625,47.109375,47.8125,48.515625,49.21875,49.921875,50.625,51.328125,52.03125,52.734375,53.4375,54.140625,54.84375,55.546875,56.25,56.953125,57.65625,58.359375,59.0625,59.765625,60.46875,61.171875,61.875,62.578125,63.28125,63.984375,64.6875,65.390625,66.09375,66.796875,67.5,68.203125,68.90625,69.609375,70.3125,71.015625,71.71875,72.421875,73.125,73.828125,74.53125,75.234375,75.9375,76.640625,77.34375,78.046875,78.75,79.453125,80.15625,80.859375,81.5625,82.265625,82.96875,83.671875,84.375,85.078125,85.78125,86.484375,87.1875,87.890625,88.59375,89.296875,90;
    lon=1.40625,2.8125,4.21875,5.625,7.03125,8.4375,9.84375,11.25,12.65625,14.0625,15.46875,16.875,18.28125,19.6875,21.09375,22.5,23.90625,25.3125,26.71875,28.125,29.53125,30.9375,32.34375,33.75,35.15625,36.5625,37.96875,39.375,40.78125,42.1875,43.59375,45,46.40625,47.8125,49.21875,50.625,52.03125,53.4375,54.84375,56.25,57.65625,59.0625,60.46875,61.875,63.28125,64.6875,66.09375,67.5,68.90625,70.3125,71.71875,73.125,74.53125,75.9375,77.34375,78.75,80.15625,81.5625,82.96875,84.375,85.78125,87.1875,88.59375,90,91.40625,92.8125,94.21875,95.625,97.03125,98.4375,99.84375,101.25,102.65625,104.0625,105.46875,106.875,108.28125,109.6875,111.09375,112.5,113.90625,115.3125,116.71875,118.125,119.53125,120.9375,122.34375,123.75,125.15625,126.5625,127.96875,129.375,130.78125,132.1875,133.59375,135,136.40625,137.8125,139.21875,140.625,142.03125,143.4375,144.84375,146.25,147.65625,149.0625,150.46875,151.875,153.28125,154.6875,156.09375,157.5,158.90625,160.3125,161.71875,163.125,164.53125,165.9375,167.34375,168.75,170.15625,171.5625,172.96875,174.375,175.78125,177.1875,178.59375,180,181.40625,182.8125,184.21875,185.625,187.03125,188.4375,189.84375,191.25,192.65625,194.0625,195.46875,196.875,198.28125,199.6875,201.09375,202.5,203.90625,205.3125,206.71875,208.125,209.53125,210.9375,212.34375,213.75,215.15625,216.5625,217.96875,219.375,220.78125,222.1875,223.59375,225,226.40625,227.8125,229.21875,230.625,232.03125,233.4375,234.84375,236.25,237.65625,239.0625,240.46875,241.875,243.28125,244.6875,246.09375,247.5,248.90625,250.3125,251.71875,253.125,254.53125,255.9375,257.34375,258.75,260.15625,261.5625,262.96875,264.375,265.78125,267.1875,268.59375,270,271.40625,272.8125,274.21875,275.625,277.03125,278.4375,279.84375,281.25,282.65625,284.0625,285.46875,286.875,288.28125,289.6875,291.09375,292.5,293.90625,295.3125,296.71875,298.125,299.53125,300.9375,302.34375,303.75,305.15625,306.5625,307.96875,309.375,310.78125,312.1875,313.59375,315,316.40625,317.8125,319.21875,320.625,322.03125,323.4375,324.84375,326.25,327.65625,329.0625,330.46875,331.875,333.28125,334.6875,336.09375,337.5,338.90625,340.3125,341.71875,343.125,344.53125,345.9375,347.34375,348.75,350.15625,351.5625,352.96875,354.375,355.78125,357.1875,358.59375,360;
    lev=1.40625,2.8125,4.21875,5.625,7.03125,8.4375,9.84375,11.25,12.65625,14.0625,15.46875,16.875,18.28125,19.6875,21.09375,22.5,23.90625,25.3125,26.71875,28.125,29.53125,30.9375,32.34375,33.75,35.15625,36.5625,37.96875,39.375,40.78125,42.1875,43.59375,45;
time=1,2,3,4,5,6,7,8;
}
