// Purpose: CDL file to generate netCDF test file

// Usage:
// ncgen -b -o in.nc in.cdl
// ncgen -b -o $HOME/nc/nco/data/in.nc $HOME/nc/nco/data/in.cdl
// mswrite -t 365 in.nc /ZENDER/tmp/in.nc
// mswrite -t 365 in.nc /ZENDER/tmp/h0001.nc
// mswrite -t 365 in.nc /ZENDER/tmp/h0002.nc
// mswrite -t 365 in.nc /ZENDER/tmp/h0003.nc
// mswrite -t 365 in.nc /ZENDER/tmp/h0004.nc
// msrcp -period 365 in.nc mss:/ZENDER/tmp/in.nc
// msrcp -period 365 in.nc mss:/ZENDER/tmp/h0001.nc
// msrcp -period 365 in.nc mss:/ZENDER/tmp/h0002.nc
// msrcp -period 365 in.nc mss:/ZENDER/tmp/h0003.nc
// msrcp -period 365 in.nc mss:/ZENDER/tmp/h0004.nc

// NB: Changing the values of the variables below, especially the coordinate 
// variables, may affect the outcome of the test script nco_tst.sh.

// NCL usage:
// id_in=addfile("/home/zender/nc/nco/data/in.nc","r")
// print(id_in)
// list_filevars(id_in)

netcdf in {
dimensions:
	band=2,lat=2,lev=3,rlev=3,lon=4,char_dim_lng=80,char_dim_sml=4,fl_dim=3,time=unlimited;
variables:
	:convention = "NCAR-CSM";
	:history = "History global attribute.\n";
	:julian_day = 200000.04;
	:RCS_Header = "$Header: /data/zender/nco_20150216/nco/data/in.cdl,v 1.15 2000-02-03 16:56:20 zender Exp $";

	float lat(lat);
	float lat_var(lat);
	float lat_wgt(lat);
	float lev(lev);
	lev:purpose = "Monotonically increasing coordinate pressure";
	float rlev(rlev);
	rlev:purpose = "Monotonically decreasing coordinate pressure";
	float lon(lon);
	double time(time);

	char fl_dim(fl_dim);
	fl_dim:long_name = "Character coordinate";
	fl_dim:units = "[chr]";

	long nbdate;
	nbdate:long_name = "base date as 6 or 8 digit integer (YYMMDD or YYYYMMDD)";
	long date(time);
	date:long_name = "current date as 6 or 8 digit integer (YYMMDD or YYYYMMDD)";

	float msk_prt_mss_prt(lon);
	msk_prt_mss_prt:long_name = "partial mask, partial missing value example";
	msk_prt_mss_prt:missing_value = 1.0e36f;

	float mss_val(lon);
	mss_val:long_name = "partial missing value example";
	mss_val:missing_value = 1.0e36f;

	float no_mss_val(lon);
	no_mss_val:long_name = "no missing value";

	float val_one_mss(lat);
	val_one_mss:long_name = "one regular value, one missing value";
	val_one_mss:missing_value = 1.0e36f;

	float wgt_one(lat);
	wgt_one:long_name = "all values are one";

	float mss_val_all(lon);
	mss_val_all:long_name = "all missing values example";
	mss_val_all:missing_value = 1.0e36f;

	float scalar_var;
	scalar_var:long_name = "scalar variable";
	scalar_var:units = "Fraction";

	float float_var;
	float_var:long_name = "float";

	double double_var;
	double_var:long_name = "double";

	long long_var;
	long_var:long_name = "long";

	short short_var;
	short_var:long_name = "short";

	char char_var;
	char_var:long_name = "char";

	char char_var_space;
	char_var_space:long_name = "Character variable with whitespace on ends";

	char char_var_nul;
	char_var_nul:long_name = "Character variable containing one NUL";

	char char_var_multinul(lev);
	char_var_multinul:long_name = "Character variable containing multiple NULs";

	char fl_nm(char_dim_lng);
	fl_nm:long_name = "Variable contains a file name";

	char fl_nm_arr(fl_dim,char_dim_lng);
	fl_nm_arr:long_name = "Variable that contains a short array of file names";
	fl_nm_arr:units = "[sng]";

	char non_nul_trm_char_one_dim(char_dim_sml);
	non_nul_trm_char_one_dim:long_name = "Variable contains a one-dimensional array of characters that is not NUL-terminated";
	non_nul_trm_char_one_dim:units = "[chr]";

	char non_nul_trm_char_two_dim(fl_dim,char_dim_sml);
	non_nul_trm_char_two_dim:long_name = "Variable contains a two-dimensional array of characters that are not NUL-terminated";
	non_nul_trm_char_two_dim:units = "[chr]";

	byte byte_var;
	byte_var:long_name = "byte";

	float zero;
	zero:long_name = "zero";

	float one;
	one:long_name = "one";

	float two;
	two:long_name = "two";

	float three;
	three:long_name = "three";

	float negative_one;
	negative_one:long_name = "negative one";

	float lev_var(lev);
	lev_var:long_name = "lev_var";

	float lev_wgt(lev);
	lev_wgt:long_name = "lev_wgt";

	float g;
	g:long_name = "g";

	float z(lev);
	z:long_name = "Height";
	z:units = "meter";
	z:purpose = "Height stored with a monotonically increasing coordinate";

	float rz(rlev);
	rz:long_name = "Height";
	rz:units = "meter";
	rz:purpose = "Height stored with a monotonically decreasing coordinate";

	float one_dim_var(band);

	float att_var;
	att_var:byte_att = '\0';
	att_var:char_att = "Sentence one.\nSentence two.\n";
	att_var:short_att = 37s;
	att_var:long_att = 73l;
	att_var:float_att = 73.0f,72.0f,71.0f;
	att_var:double_att = 73.0d;

	long band_var(lev,band);
	band_var:byte_att = '\0';
	band_var:char_att = "Sentence one.\nSentence two.\n";
	band_var:short_att = 37s;
	band_var:long_att = 73l;
	band_var:float_att = 73.f;
	band_var:double_att = 73.d;

	float three_dim_var(lat,lev,lon);
	three_dim_var:long_name = "three dimensional variable";
	three_dim_var:units = "Fraction";

	float two_dim_var(lat,lev);
	two_dim_var:long_name = "two dimensional variable";
	two_dim_var:units = "Fraction";

	float mask(lat,lon);
	mask:long_name = "mask variable like ORO";
	mask:units = "Fraction";

	float ORO(lat,lon);
	ORO:long_name = "Orography";
	ORO:units = "Fraction";

	float weight(lat);
	weight:long_name = "Gaussian weight";
	weight:units = "Fraction";

	float gw(lat);
	gw:long_name = "gw variable like gw";
	gw:units = "Fraction";

	float rec_var_flt(time);
	rec_var_flt:long_name = "record variable, float";

	double rec_var_dbl(time);
	rec_var_dbl:long_name = "record variable, double";

	long one_dim_rec_var(time);
	one_dim_rec_var:long_name = "one dimensional record variable";
	one_dim_rec_var:units = "second";

	float tpt(time);
	tpt:long_name = "one dimensional record variable";
	tpt:units = "second";

	float rec_var_flt_mss_val_flt(time);
	rec_var_flt_mss_val_flt:long_name = "record variable, float, with float missing values";
	rec_var_flt_mss_val_flt:missing_value = 1.0e36f;

	float rec_var_flt_mss_val_dbl(time);
	rec_var_flt_mss_val_dbl:long_name = "record variable, float, with double missing values";
	rec_var_flt_mss_val_dbl:missing_value = 1.0e36d;

	char one_dim_rec_var_sng(time);
	one_dim_rec_var_sng:long_name = "one dimensional record variable of string";

	float time_lon(time,lon);
	time_lon:long_name = "Record variable of longitude coordinate";

	char two_dim_rec_var_sng(time,lev);
	two_dim_rec_var_sng:long_name = "two dimensional record variable of string";

	float two_dim_rec_var(time,lev);
	two_dim_rec_var:long_name = "two dimensional record variable";
	two_dim_rec_var:units = "watt meter-2";

	float three_dim_rec_var(time,lat,lon);
	three_dim_rec_var:long_name = "three dimensional record variable";
	three_dim_rec_var:units = "watt meter-2";

	float four_dim_rec_var(time,lat,lev,lon);
	four_dim_rec_var:long_name = "four dimensional record variable";
	four_dim_rec_var:units = "watt meter-2";

data:
	ORO=1.,1.,1.,1.,1.,1.,1.,1.;
	att_var=10.;
	band_var=1,2,3,4,5,6;
	byte_var='z';
	char_var="z";
	char_var_space=" ";
	char_var_nul='\0';
	char_var_multinul="\b\n\0";
	double_var=10.;
	fl_nm="/home/zender/nc/nco/data/in.cdl";
	fl_dim="a","b","3";
	float_var=10.;
	g=9.8;
	gw=10.,10.;
	lat=-90,90;
	lat_var=1.,2.;
	lat_wgt=1.,2.;
	lev=100,500,1000;
	lev_var=100.,500.,1000.;
	lev_wgt=10,2,1;
	lon=0,90,180,270;
	mask=0.,1.,0.,0.,1.,1.,0.,2.;
//	mask=0.,0.,0.,0.,0.,0.,0.,0.;
//	mask=1.,1.,1.,1.,1.,1.,1.,1.;
	msk_prt_mss_prt=0.5,1.0e36,1.5,1.0e36;
	mss_val=73,1.0e36,73,1.0e36;
	mss_val_all=1.0e36,1.0e36,1.0e36,1.0e36;
	negative_one=-1.;
	no_mss_val=73,1.0e36,73,1.0e36;
	non_nul_trm_char_one_dim='a','b';
	non_nul_trm_char_two_dim="abcd","efgh","ijkm";
	one=1.;
	one_dim_rec_var=1,2,3,4,5,6,7,8,9,10;
	tpt=273.1,273.2,273.3,273.4,273.5,273.6,273.7,273.8,273.9,273.10;
	one_dim_rec_var_sng="Hello Wor";
	one_dim_var=1.,10.;
	rec_var_dbl=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	rec_var_flt=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	rec_var_flt_mss_val_dbl=1.0e36,2.,3.,4.,5.,6.,7.,8.,1.0e36,1.0e36;
	rec_var_flt_mss_val_flt=1.0e36,2.,3.,4.,5.,6.,7.,8.,1.0e36,1.0e36;
	rlev=1000,500,100;
	rz=0,5000,17000;
	scalar_var=10.;
	short_var=10;
	three=3.;
	three_dim_var=0.,1.,2.,3.,4.,5.,6.,7.,8.,9.,10.,11.,12.,13.,14.,15.,16.,17.,18.,19.,20.,21.,22.,23.;
	time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	two=2.;
	two_dim_var=1.5,5.5,9.5,13.5,17.5,21.5;
	val_one_mss=1.,1.0e36;
	weight=10.,10.;
	wgt_one=1.,1.;
	z=17000,5000,0;
	zero=0.;
 	date=640312,640313,640314,640315,640316,640317,640318,640319,640320,640321;
 	long_var=10;
 	nbdate=640312;
	fl_nm_arr="/data/zender/dstccm04/dstccm04_8589_01.nc",
		"/data/zender/dstccm04/dstccm04_8589_02.nc",
		"/data/zender/dstccm04/dstccm04_8589_03.nc";
	time_lon=0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0,
			0.0,90.0,180.0,270.0;
	two_dim_rec_var_sng="abc",
				"bcd",
				"cde",
				"def",
				"efg",
				"fgh",
				"ghi",
				"hij",
				"jkl",
				"klm";
	two_dim_rec_var=1.,2.0,3.,
			1.,2.1,3.,
			1.,2.2,3.,
			1.,2.3,3.,
			1.,2.4,3.,
			1.,2.5,3.,
			1.,2.6,3.,
			1.,2.7,3.,
			1.,2.8,3.,
			1.,2.9,3.;
	three_dim_rec_var= 	 1, 2, 3, 4, 5, 6, 7, 8,
				 9,10,11,12,13,14,15,16,
				17,18,19,20,21,22,23,24,
				25,26,27,28,29,30,31,32,
				33,34,35,36,37,38,39,40,
				41,42,43,44,45,46,47,48,
				49,50,51,52,53,54,55,56,
				57,58,59,60,61,62,63,64,
				65,66,67,68,69,70,71,72,
				73,74,75,76,77,78,79,80;
	four_dim_rec_var= 	  1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12,
				 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24,
				 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36,
				 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48,
				 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60,
				 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72,
				 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84,
				 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96,
				 97, 98, 99,100,101,102,103,104,105,106,107,108,
				109,110,111,112,113,114,115,116,117,118,119,120,
				121,122,123,124,125,126,127,128,129,130,131,132,
				133,134,135,136,137,138,139,140,141,142,143,144,
				145,146,147,148,149,150,151,152,153,154,155,156,
				157,158,159,160,161,162,163,164,165,166,167,168,
				169,170,171,172,173,174,175,176,177,178,179,180,
				181,182,183,184,185,186,187,188,189,190,191,192,
				193,194,195,196,197,198,199,200,201,202,203,204,
				205,206,207,208,209,210,211,212,213,214,215,216,
				217,218,219,220,221,222,223,224,225,226,227,228,
				229,230,231,232,233,234,235,236,237,238,239,240;
}

