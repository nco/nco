�HDF

         ����������     0       .��OHDRx"     P      �      z      �      
         �      G       )         _nc3_strict                '        Conventions          CF-1.0$       history         Fri Jan 16 16:52:29 2015: ncks -O -7 --cnk_dmn time,10 in_4c.nc in.cdl
Tue Jan 13 13:29:14 2015: ncks -O -7 --cnk_dmn time,10 ../data/in.nc ../data/in_4c.nc
History global attribute.
Attributes like this often have embedded newlines to enhance legibility.
Such newlines should serve as linebreaks on the screen, hence,
friendly CDL converters print a single NC_CHAR attribute as a comma-separated list of strings
where each embedded delimiter marks a linebreak.
Otherwise it would be harder for humans to read the CDL. D        julian_day  ?      @ 4 4�                ��Q jA(        RCS_Header          $Header: /data/zender/nco_20150216/nco/data/in.cdl,v 1.203 2015-01-17 00:53:13 zender Exp $"        NCO    	      20150117            N!OHDR                        
   *     �|   ؈             �                                                                                                                                                                                  ���OCHK     ������������������������                            �l�OHDR                        
   *     �|   ܈             �                                                                                                                                                                                  �'��OCHK+        _Netcdf4Dimid                �b)        OHDR                        
   *     �|   ��             �                                                                                                                                                                                  �7IBTHD       d(_�              q�t                             OHDR                        
   *     �|   �             �                                                                                                                                                                                  gfOCHK+        _Netcdf4Dimid                3�pw           OHDR                        
   *     �|   �             �                                                                                                                                                                                  f�OCHK+        _Netcdf4Dimid                I��F           OHDR                        
   *     �|   �             �                                                                                                                                                                                  H�c�OCHK(        units          degrees_northV�e�            OHDR                       ?      @ 4 4�     *         �G    D�     �            ������������������������+         CLASS          DIMENSION_SCALE         NAME          Lat     �                                �
aqOCHK+        _Netcdf4Dimid             
   �'z       OCHK+        _Netcdf4Dimid                 '    
    long_name          Latitude(        units          degrees_northh        purpose    K      Latitude paired with Longitude coordinate originally stored as -180 to 180.�޹gOHDR $                                    ?      @ 4 4�     *         �G    .      �            ������������������������Z     
    long_name    ;      2D variable originally stored on -180 to 180 longitude grid 
              FB,xBTHD 	      d(_�              =F4�                             OCHK    ��     �       #        units          fraction_        purpose    B      Demonstrate remapping of [-180,180) to [0,360) longitude-grid data  ���hOHDR                       ?      @ 4 4�     *         �G          ,           ������������������������+         CLASS          DIMENSION_SCALE         NAME          Lon           9                           +r��FRHP               ��������      �       @       (       (      P                                                        �G      �s�BTHD      d(-B       P      a� �BTHD      d(�1      	 P      *���FSHD  Y                             P x          �o     m       m       X�V>BTLF C�   �   /�=  �  # bO# �   zn �   �7� �   h]E e  & �j� �    E�3 B    %�� �$  ! �? `   �. 2   ߋ< �   "�~ 8   �,% �   �| c   ʊ� e  1 *�� 0   v�;	 R   h�� }#   �1�     vq� �    �� �   �̻ '   g@� �   L� �   �� =   �?6 �   SČ   # *�� �  " ��� y   Xb� �   =�� �#   ��� �    L� �    }& v   h0� V   �58 �  0 ٠�   -  !E o  6 ��H +   Y� �!   V�% �$   �| y  * N�J                             BTLF                      ,            B            [            u            �            �            �            �    	        �    
                              ,           @           V           m           �           �           �           �           �                      +           A           V           l           �           �           �           �           �           �               +XI�       OCHK    ��     �       (    
    long_name    	      Longitude"        units          degreesR        purpose    5      Longitude coordinate originally stored as -180 to 180X        notes    =      Longitude = [-180.0,180.0) is not CF-compliant, yet is common  \��OHDR*$                                                
   *     �|    h�     �            ������������������������m     
    long_name    N      Orography, an enumerated yet continuous type: ocean=0.0, land=1.0, sea ice=2.0#        units          fraction  (% OHDR                        
   *     �|   ��                 ������������������������1     
    long_name          reference pressure!        units          pascal .                                                  +Q4pOHDR4    
                     ��������                  �     �       
   +     �|   ؐ     
                 ������������������������/     
    long_name          surface pressure!        units          pascal    �7}�OHDR                        
   *     �|   ��             �                                                                                                                                                                                  �B�OHDR                        
   *     �|   ��             �                                                                                                                                                                                  ���OHDR                        
   *     �|   ��             �                                                                                                                                                                                  } YOHDR                        
   *     �|   ��             �                                                                                                                                                                                  �� OHDR                        
   *     �|   ��             �                                                                                                                                                                                  VK��OHDR                        
   *     �|   ��             �                                                                                                                                                                                  8��OHDR                        
   *     �|   ��             �                                                                                                                                                                                  ��`�OHDR                        
   *     �|   ��             �                                                                                                                                                                                  _Z��OHDR                        
   *     �|   ��             �                                                                                                                                                                                  �Æ�OHDR                        
   *     �|   ��             �                                                                                                                                                                                  �p�LOHDR                        
   *     �|   ��             �                                                                                                                                                                                  �vuOHDR                        
   *     �|   ��             �                                                                                                                                                                                  -p�OHDR                        
   *     �|   ��             �                                                                                                                                                                                  �]!XOHDR                        
   *     �|   ��             �                                                                                                                                                                                  ��OHDR                        
   *     �|   ��             �                                                                                                                                                                                  _�eOHDR                        
   *     �|   ��             �                                                                                                                                                                                  �RVOHDR                        
   *     �|   ĉ             �                                                                                                                                                                                  ��LOHDR                        
   *     �|   ȉ             �                                                                                                                                                                                  Bc xOHDR                        
   *     �|   ̉             �                                                                                                                                                                                  N��OHDR                        
   *     �|   Љ             �                                                                                                                                                                                  )>P+OHDR                        
   *     �|   ԉ             �                                                                                                                                                                                  ;��hOHDR                        
   *     �|   ؉             �                                                                                                                                                                                  �?�7BTIN !           C        A   e        I	   �        �  # �        �   �        J   �        �  .        �   /       �!         !�3      !5]      !̈́      !�      !��      !�     !5C     !�     �      �o`     m           �           �           �           �           �                      +           A           V           l           �           �           �           �           �           �               +XI�       BTLF "        3   #        I   $        _   %        u   &        �   '        �   (        �   )        �   *        �   +           ,        +   -        A   .        W   /        m   0        �   1        �   2        �   3        �   4        �   5        �   6           7           8        3   9        I   :        _   ;        u   <        �   =        �   >        �   ?        �   @        �   A           B        +   k��       OHDR                        
   *     �|   ܉             �                                                                                                                                                                                  ��(�OHDR                        
   *     �|   ��             �                                                                                                                                                                                  N��OHDR                        
   *     �|   �             �                                                                                                                                                                                  ���jOHDR                        
   *     �|   �             �                                                                                                                                                                                  �m[�OHDR                        
   *     �|   �             �                                                                                                                                                                                  ��ϺOHDR                        
   *     �|   ��             �                                                                                                                                                                                  [s#�OHDR                        
   *     �|   �             �                                                                                                                                                                                  �t�OHDR                        
   *     �|   ��             �                                                                                                                                                                                  ��jOHDR                        
   *     �|   ��             �                                                                                                                                                                                  �5s�OHDR                        
   *     �|    �             �                                                                                                                                                                                  �6#OHDR                        
   *     �|   �             �                                                                                                                                                                                  #�Q
OHDR                        
   *     �|   �             �                                                                                                                                                                                  ��N�BTIN ���  �    8�>    C�`b .  2 ���z ?  & ���� �   j6]�    �� A         +1&     +�      +�     +-D      +Ux      ,�      -7r     ?r2 �| c   ʊ� e  1 *�� 0   v�;	 R   h�� }#   �1�     vq� �    �� �   �̻ '   g@� �   L� �   �� =   �?6 �   SČ   # *�� �  " ��� y   Xb� �   =�� �#   ��� �    L� �    }& v   h0� V   �58 �  0 ٠�   -  !E o  6 ��H +   Y� �!   V�% �$   �| y  * N�J                             BTLF �׊| �   qoD} T   ��~ �   �Q�� y    QO� 3   9Y � �#   [�ׄ �
   %z�� �"  " !Q� �   eL�� �   )� �   PG4� �   �Tl� I	   �Yt� �   [)� C   ��9�    �f�� �   �`É �   g�&�   * �W� :!   �،� �"   n�΍ �   Ͱݍ t   �M� �   U�)� �   ~�*� �   �ˑ I   A�ȓ A   �Eܓ v   mʔ m   ��A� m   pXe�     ��    �yE� m!   ��ӗ �   5��    �t�� #   ���� !  & �_�� p   fE*�    E�$� �   `�o� m   �b� �  &  ��U                             OHDR                        
   *     �|   �             �                                                                                                                                                                                  � ��OHDR                        
   *     �|   �             �                                                                                                                                                                                   N&OHDR                        
   *     �|   �             �                                                                                                                                                                                  ��$�OHDR                        
   *     �|   �             �                                                                                                                                                                                  7�,�OHDR                        
   *     �|   �             �                                                                                                                                                                                  T��OHDR                        
   *     �|    �             �                                                                                                                                                                                  ��]�OHDR                        
   *     �|   $�             �                                                                                                                                                                                  Gq�hOHDR                        
   *     �|   (�             �                                                                                                                                                                                  ��~,OHDR                        
   *     �|   ,�             �                                                                                                                                                                                  �v
OHDR                        
   *     �|   0�             �                                                                                                                                                                                  ��gzOHDR                        
   *     �|   4�             �                                                                                                                                                                                  �F_�OHDR                        
   *     �|   8�             �                                                                                                                                                                                  �]{kOHDR                        
   *     �|   <�             �                                                                                                                                                                                  <�F�OHDR                        
   *     �|   @�             �                                                                                                                                                                                  �l�POHDR                        
   *     �|   D�             �                                                                                                                                                                                  �/W`OHDR                        
   *     �|   H�             �                                                                                                                                                                                  AD��OHDR                        
   *     �|   L�             �                                                                                                                                                                                  ���OHDR                        
   *     �|   P�             �                                                                                                                                                                                  ����OHDR                        
   *     �|   T�             �                                                                                                                                                                                  �aOHDR                        
   *     �|   X�             �                                                                                                                                                                                  U�I�OHDR                        
   *     �|   \�             �                                                                                                                                                                                  _r��OHDR                        
   *     �|   `�             �                                                                                                                                                                                  ��BTLF D        W   E        m   F        �   G        �   H        �   I        �   J        �   K        �   L           M           N        3   O        I   P        _   Q        u   R        �   S        �   T        �   U        �   V        �   W           X        +   Y        A   Z        W   [        m   \        �   ]        �   ^        �   _        �   `        �   a        �   b        	   c        	   d        3	   �E�!       OHDR                        
   *     �|   d�             �                                                                                                                                                                                  Y��OHDR                        
   *     �|   h�             �                                                                                                                                                                                  �ݰFOHDR                        
   *     �|   l�             �                                                                                                                                                                                  �w5LOHDR                        
   *     �|   p�             �                                                                                                                                                                                  ��?OHDR                        
   *     �|   t�             �                                                                                                                                                                                  �/S9OHDR                        
   *     �|   x�             �                                                                                                                                                                                  �e&ZOHDR                        
   *     �|   |�             �                                                                                                                                                                                  �W�OHDR                        
   *     �|   ��             �                                                                                                                                                                                  '� �OHDR                        
   *     �|   ��             �                                                                                                                                                                                  ��H#OHDR                        
   *     �|   ��             �                                                                                                                                                                                  Y��^OHDR                        
   *     �|   ��             �                                                                                                                                                                                  �.jOHDR                        
   *     �|   ��             �                                                                                                                                                                                  �p]OHDR                        
   *     �|   ��             �                                                                                                                                                                                  n���OHDR                        
   *     �|   ��             �                                                                                                                                                                                  �*�uOHDR                        
   *     �|   ��             �                                                                                                                                                                                  VO��OHDR                        
   *     �|   ��             �                                                                                                                                                                                  �F�gOHDR                        
   *     �|   ��             �                                                                                                                                                                                  ڟC@OHDR                        
   *     �|   ��             �                                                                                                                                                                                  KopOHDR                        
   *     �|   ��             �                                                                                                                                                                                  ��K�OHDR                        
   *     �|   ��             �                                                                                                                                                                                  ��ϲOHDR                        
   *     �|   ��             �                                                                                                                                                                                  �	7�OHDR                        
   *     �|   ��             �                                                                                                                                                                                  �wD'OHDR                        
   *     �|   ��             �                                                                                                                                                                                  �#<fOHDR                        
   *     �|   ��             �                                                                                                                                                                                  �.BTLF �V-�    �pD� �   R*� �   <+5�    +'N� �    �2� �   " m�&� ,    ��� ^   �[��    �� W   �hw� �   ��� �    �ܶ� B   �sx� [   0Ή� �!   �έ A   �A� I   [{�� +   ��G� �  * �C� �   {3p� z   �d� C$   �� �!    �$ʹ �   i��� M"  " \��� _   �� � �!   e� �   �z� �   �/� k   K�>� %  * �Č� �   S�� l   A[�� [    ��� �	   Uy� �   �� �   ���    ��� $   �.=� �    T�� �   �Z�� 	   �L� �   Z�� u	   ����                  OHDR                        
   *     �|   Ċ             �                                                                                                                                                                                  ��r�OHDR                        
   *     �|   Ȋ             �                                                                                                                                                                                  ��+�OHDR                        
   *     �|   ̊             �                                                                                                                                                                                  v�"OHDR                        
   *     �|   Њ             �                                                                                                                                                                                  �'<OHDR                        
   *     �|   Ԋ             �                                                                                                                                                                                  u �OHDR                        
   *     �|   ؊             �                                                                                                                                                                                  ���OHDR                        
   *     �|   ܊             �                                                                                                                                                                                  ��NgOHDR                        
   *     �|   ��             �                                                                                                                                                                                  ˷XOHDR                        
   *     �|   �             �                                                                                                                                                                                  v~��OHDR                        
   *     �|   �             �                                                                                                                                                                                  *~BTLF f        _	   g        u	   h        �	   i        �	   j        �	   k        �	   l        �	   m        
   n        +
   o        A
   p        W
   q        m
   r        �
   s        �
   t        �
   u        �
   v        �
   w        �
   x           y        '   z        A   {        [   |        t   }        �   ~        �           �   �        �   �           �        0   �        O  ! �        p   �        �   �        �  # O�T>       OHDR                        
   *     �|   �             �                                                                                                                                                                                  ��6iOHDR                        
   *     �|   ��             �                                                                                                                                                                                  ��i(OHDR                        
   *     �|   �             �                                                                                                                                                                                  x�pOHDR                        
   *     �|   ��             �                                                                                                                                                                                  Pj�GOHDR                        
   *     �|   ��             �                                                                                                                                                                                  [&OHDR                        
   *     �|    �             �                                                                                                                                                                                  ��UYOHDR                        
   *     �|   �             �                                                                                                                                                                                  X&N�OHDR                        
   *     �|   �             �                                                                                                                                                                                  =��OHDR                        
   *     �|   �             �                                                                                                                                                                                  R��OHDR                        
   *     �|   �             �                                                                                                                                                                                  n��OHDR                        
   *     �|   �             �                                                                                                                                                                                  L�	OHDR                        
   *     �|   �             �                                                                                                                                                                                  ��%6OHDR                        
   *     �|   �             �                                                                                                                                                                                  �eOHDR                        
   *     �|    �             �                                                                                                                                                                                  rܐ�OHDR                        
   *     �|   $�             �                                                                                                                                                                                  $���OHDR     
       ��������            
   +     �   �     
           ������������������������L         DIMENSION_LIST                              D�        +        _Netcdf4Dimid                      �(�OHDR                                   
   *     �|   (�                 ������������������������#     
    long_name          area!        units          meter2    k�     Z           |     9             5��7OHDR                                   
   *     �|    �A     Q            ������������������������-     
    long_name          area version 2!        units          meter2    ��     Z                          있JOHDR                                   
   *     �|    �A     Q            ������������������������.     
    long_name          area asymmetric!        units          meter2    d�     Z                         i#nOHDR�    
       ��������                
   +     �|    	 V     �
     �!        H�     
          ��������
                                                :                                                             5                                                        5                                                        6                                                         W                                                                                          t                                                                                                                       �|�OHDR@$                                            
   *     �    	 ��     ��     4�        @�             �   ��������                                          :                                                             5                                                        5                                                        6                                                         ?                                                                  D                                                                       O� �OHDR $                                              *   �   X�                 ������������������������\         DIMENSION_LIST                              D�           D�            �	      9            cc�mOHDR 4                                                            *   �   `�                 ������������������������    ��     z       +        _Netcdf4Dimid                                                      �ܔvOHDR 4    
                     ��������                            +   �   x�     
                 ������������������������    R�     z       +        _Netcdf4Dimid                                            �Y��OHDR $                                              *   �   x�                 ������������������������)     
    long_name    
      byte array    ��     j       +        _Netcdf4Dimid                      ��D�OHDR                      *   �   ��                 ������������������������#     
    long_name          byte n                                                                                                                  ����OHDR                      *   �   ��                 ������������������������,     
    long_name          negative byte e                                                                                                         �Ȯ�OHDR                    *       ��                 ������������������������#     
    long_name          char r                                                                                                                      ���OHDR                    *       ��                 ������������������������D     
    long_name    %      Character variable containing one NUL Q                                                                                     X��OHDR                    *       ��                 ������������������������I     
    long_name    *      Character variable with whitespace on ends L                                                                                �%.OHDR�                                  
   *     �|    ��     r            ������������������������>     
    long_name          test CF coordinates conventions1        coordinates          lat_gds lon_gds �        reason          Test whether coordinates attribute strings that end with a space break after nco_var_lst_crd_ass_add() call to nco_lst_prs_2d()  U��OHDR�    
       ��������                
   +     �|    ��     s            ������������������������E     
    long_name    &      test CF ancillary_variables convention4        standard_name          specific_humidityJ        ancillary_variables    !      cnv_CF_ncl_var_1 cnv_CF_ncl_var_2s        purpose    V      Main variable that has ancillary variables named cnv_CF_ncl_var_1 and cnv_CF_ncl_var_2   ��{�OHDR�    
       ��������                
   +     �|    ��     �            ������������������������E     
    long_name    &      test CF ancillary_variables conventionC        standard_name           specific_humidity standard_errorm        purpose    P      Ancillary variable for cnv_CF_ncl. Other ancillary variable is cnv_CF_ncl_var_2.   �P�]OHDR     
       ��������                
   +     �|    p=     R            ������������������������E     
    long_name    &      test CF ancillary_variables convention    �      �           ��     Z                   �J�BTLF �        �   �           �        "   �        =   �        S   �        m   �        �   �        �   �        �   �        �   �           �        -   �        E   �        ^   �        v   �        �   �        �   �        �  " �        �   �           �          # �        @   �        T   �        p   �        �   �        �   �        �   �        �   �           �        ,   �        C   �        Z   �        t   u�P       OCHKD        standard_name    !      specific_humidity detection_limitm        purpose    P      Ancillary variable for cnv_CF_ncl. Other ancillary variable is cnv_CF_ncl_var_1.�O�8OHDR     
       ��������            
   +     �    �=     R            ������������������������Y     
    long_name    :      current date as 6- or 8-digit integer (YYMMDD or YYYYMMDD)    �     Z                             �N�BTLF ���� �  $ R|+� F#   �=�� m   Z�� �  + S�� t$  ! ��� �   US�� @   ��� u   A�)� �   ��A� z   ���� �   �DT� �   ��e� :   ꫍� �  " B�� \   v�� �   k_�� �  " `��� �   i��� �   Ҭ�� �    {a�� +
   1�� �   �$�    ��� �    ��M�    . b1w� .    sE�� u    i��� �   �D� +   6W4� -   �߽� �   ���� �
   Gܗ� �  0 ��� �   .��� 0   '�;� m  6 )oM� 	   p�~� F   E>�� A   k-�    �%��    ���� S   D�� �	   �,�� �	   �)� W   ���       OHDR                               
   *     �   ��                 ������������������������H     
    long_name    )      Date (as array of ints: YYYY,MM,DD,HH,MM)    `�     Z           �W     9        
              >�9OHDR $    
              ��������                   +        ��     �                  ������������������������@     
    long_name    !      A record variable of date strings         units          [sng] 
              ���OHDR                                   
   *     �|   (     �            ������������������������+         CLASS          DIMENSION_SCALE         NAME          dgn     �      9           �      j          h�[BTLF ��? �  . :9�@ �   �s-A �   ��sA    ��B l   �@�B �  * ��B    ��C L   �QC �   � �D �   �W�D    >��E )#   Ә�F f   ��G c#   `4H    n2YI �   ){I �   n�J   * �G�K _	   K8�K D  + �L    �S~L �   1��L �   oiM (  + ��zN "   �ZO   & ��\P �  6 �8@Q    ��Q I   �g<R �#   ��LR u   CTR ,$   E�QT �  $ ~�U `    �f�W A
   Ќ|Y �   L5�Y �  2 Gd"Z �   l�s[ W   ���[ "   �Q] �   c�_ �   ;ƙ` �!   ,��E �	   �)� W   ���       OCHK\    
    long_name    =      degenerate coordinate (dgn means degenerate, i.e., of size 1)���OHDR                                   
   *     �|    j>     Q            ������������������������Z     
    long_name    ;      degenerate variable (dgn means degenerate, i.e., of size 1)    ��     Z                    �� :OHDR            ?      @ 4 4�     *         �G   ��                 ������������������������%     
    long_name          double ]                                                                                                 �� OHDR            ?      @ 4 4�     *         �G   ɋ                 ������������������������%     
    long_name          doubleD        _FillValue  ?      @ 4 4�                � y��hG                        Ԧ�_OHDR                        
   *     �|   ы                 ������������������������-     
    long_name          Dry Deposition Y                                                                                             6m�OHDR                        
   *     �|   Ջ                 ������������������������/     
    long_name          Total Deposition W                                                                                           D���OHDR                        
   *     �|   ً                 ������������������������-     
    long_name          Wet Deposition Y                                                                                             �ga�OHDR            ?      @ 4 4�     *         �G   ݋                 ������������������������8     
    long_name          e, natural logarithm base J                                                                              2W�OCHK+        _Netcdf4Dimid                ��~                    OHDR                        
   *     �|   �                 ������������������������8     
    long_name          e, natural logarithm base N                                                                                  ��:LOHDRW                              *       *     �            ������������������������+         CLASS          DIMENSION_SCALE !        NAME          fl_dmn +        _Netcdf4Dimid                3    
    long_name          Character coordinate         units          [chr]  .OHDR     P       P                   *       �     P            ������������������������<     
    long_name          Variable contains a file name    �     Z       +        _Netcdf4Dimid                       �i�OHDR $           P              P                   *        ��     �            ������������������������Q     
    long_name    2      Variable that contains a short array of file names         units          [sng]      ���OHDR $    
       P       ��������P                   +        ^�     �                  ������������������������>     
    long_name          A record variable of file names         units          [sng]                 �_|OHDR                                   
   *     �|    �     r            ������������������������1     
    long_name          _FillValue example@        _FillValue                             �y�      e$g�OHDRD                                  
   *     �|    ��     r            ������������������������1     
    long_name          _FillValue example@        _FillValue                             �y�C        missing_value                             �y�  ���_OHDR                        
   *     �|   L�                 ������������������������$     
    long_name          float b                                                                                                      ��f�OHDR                        
   *     �|   P�                 ������������������������#     
    long_name          four c                                                                                                       /�Z�OHDR-D    
                            ��������                         `�     �       
   +     �|   ��     
                    ������������������������?     
    long_name           four dimensional record variable'        units          watt meter-2    �� �OHDR                        
   *     �|   T�                 ������������������������      
    long_name          g f                                                                                                          �N�XOHDR�$    
              ��������           M�     �       
   +     �|   0�     
              ������������������������0     
    long_name          Geodesic variable         units          meter0        coordinates          lat_gds lon_gds]        purpose    @      Test auxiliary coordinates like those that define geodesic grids    �}]EOHDR                                  
   *     �|  
 Q     �            ������������������������+         CLASS          DIMENSION_SCALE "        NAME          gds_crd +        _Netcdf4Dimid                2    
    long_name          Geodesic coordinate!        units          degreei        purpose    L      enumerated coordinate like those that might define points in a geodesic grid0        coordinates          lat_gds lon_gds  ΢l�OHDRs                                  
   *     �|    �     r            ������������������������0     
    long_name          Geodesic variable         units          meter]        purpose    @      Test auxiliary coordinates like those that define geodesic grids0        coordinates          lat_gds lon_gds  �绵OHDR�                                  
   *     �|    ��     r            ������������������������G     
    long_name    (      Geodesic variable on non-coordinate grid         units          meter�        purpose    }      Test auxiliary coordinates like those that define geodesic grids but where underlying dimension is a non-coordinate dimension8        coordinates          lat_gds_ncd lon_gds_ncd   �(�OHDR                                   
   *     �|    �@     Q            ������������������������2     
    long_name          gw variable like gw#        units          fraction    �     Z                   :2OOHDR     @       @                       
   *     �|    JA     Q            ������������������������6     
    long_name          gw variable like gw_T42#        units          fraction    (�     Z               ��]OHDR                                   
   *     �|   ��                 ������������������������F     
    long_name    '      hybrid A coefficient at layer midpoints    ��     Z           ��      9                �?pOCHKB        scale_factor                              �?���;      OHDR                                   
   *     �|   ̎                 ������������������������F     
    long_name    '      hybrid B coefficient at layer midpoints    �     Z           �A     9                (�OHDR $                                                
   *     �|   ؎                 ������������������������?         purpose    "      Cell boundaries for lev coordinate    m�     j           �A     9        olhOHDR                    
   *     �   ��                 ������������������������"     
    long_name          int l                                                                                                                Ƃ��OHDR�                                  
   *     �|  1 �I     R          3 ������������������������+         CLASS          DIMENSION_SCALE         NAME          lat +        _Netcdf4Dimid                =    
    long_name          Latitude (typically midpoints)(        units          degrees_north#        bounds          lat_bnd  �FM�OHDR                                   
   *     �|    i      r            ������������������������S     
    long_name    4      Latitude for 2D rectangular grid stored as 1D arrays    O      6                           �u�MBTLF �        �   �        �   �        �   �        �   �           �        2   �        L   �        f   �        �   �        �   �        �    �        �  $ �        �   �           �        0   �        F   �        `   �        z   �        �   �        �   �        �   �        �   �           �           �        8   �        R   �        l   �        �   �        �   �        �   �        �   �           �        0   ��B       OHDR                                  
   *     �|    m     r            ������������������������Q     
    long_name    2      Latitude for 2D irregular grid stored as 1D arrays(        units          degrees_north  ݂}OHDR$                                                
   *     �|    �      �            ������������������������R     
    long_name    3      Latitude for 2D rectangular grid stored as 2D array(        units          degrees_north  ,��
OHDR$                                                
   *     �|    ;�     �            ������������������������P     
    long_name    1      Latitude for 2D irregular grid stored as 2D array(        units          degrees_north  �Q�HOHDR    @       @                       
   *     �|    ��     �            ������������������������+         CLASS          DIMENSION_SCALE "        NAME          lat_T42 +        _Netcdf4Dimid                  �إ�OHDR $                                                
   *     �|   |�                 ������������������������?         purpose    "      Cell boundaries for lat coordinate    ��     j           QC     9        �3��OHDR�    
       
           ?      @ 4 4�     *         �G   h     P            ������������������������+         CLASS          DIMENSION_SCALE "        NAME          lat_cal +        _Netcdf4Dimid                &    
    long_name          lat_cal/        units          days since 1964-2-28%    	    calendar          360_day�qW�OHDR                                   
   *     �|   ��                 ������������������������L         DIMENSION_LIST                              D�     [       �C     9                                {�f_OHDRh                      ?      @ 4 4�     *         �G    ��     r            ������������������������'     
    long_name          Latitude+        standard_name          latitude!        units          degree[        purpose    >      1-D latitude coordinate referred to by geodesic grid variables  �K�bOHDR                      ?      @ 4 4�     *         �G    C     r            ������������������������'     
    long_name          Latitude+        standard_name          latitude!        units          degreer        purpose    U      1-D latitude coordinate referred to by "non-coordinate" (ncd) geodesic grid variables  �H�OHDR                                  
   *     �|   �                 ������������������������+         CLASS          DIMENSION_SCALE "        NAME          lat_grd +        _Netcdf4Dimid                C    
    long_name    $      Latitude grid (typically interfaces)(        units          degrees_north�v��OHDR�                              
   *     �   �     �           
 ������������������������+         CLASS          DIMENSION_SCALE (        NAME          lat_times_lon +        _Netcdf4Dimid                v    
    long_name    W      Element index (i.e., C-based storage order) for 2D coordinate grids stored as 1D arrays  �H��OHDR[                   
   *     �   Ԑ                 �������������������������     
    long_name    �      Number of elements in 2D coordinate grids. Rectangular and irregular test grids have this many total elements. The coordinates and elements are stored as 1D or 2D arrays for grid types 1D and 2D respectively.PR�xOHDR                                   
   *     �|   $                 ������������������������L         DIMENSION_LIST                              D�     ^       eD     9                                �ڶkOHDR                                   
   *     �|   ,                 ������������������������L         DIMENSION_LIST                              D�     _       �D     9                                �љ�OHDR�                                  
   *     �|   4                 {�      `      �       w                                                                                                                                                                                                                                                                                                                                                                                          �Q��FRHP               ���������       �                                                                                  (  �t       ���pFSHD  �                              P x (        Ś                   G��"BTLF  %        ���     +      ��< �      
   2�y A         _��� D        yHT� _    +     e>� �    I     o�E� �    0      i�� �   |    �� �     	   �U��    "     �!� c        �����%�                                                                                                                                                                                                                                                                                                          BTLF 	     +       A          _    +      �    I      �    0         "      %         D         c         �     	    �      
    �   |    {'�                                                                                                                                                                                                                                                                                                                                                          OHDR                                   
   *     �|   @                 ������������������������L         DIMENSION_LIST                              D�     `       �D     9                                ��_OHDR                                   
   *     �|    E     Q            ������������������������&     
    long_name          lev_varL        DIMENSION_LIST                              D�     a         S%�hOHDR                                   
   *     �|    aE     Q            ������������������������&     
    long_name          lev_wgtL        DIMENSION_LIST                              D�     b         ��OHDRu                                  
   *     �|  + M               - ������������������������+         CLASS          DIMENSION_SCALE         NAME          lon +        _Netcdf4Dimid                >    
    long_name          Longitude (typically midpoints)'        units          degrees_east  �"�OHDR                                  
   *     �|    ��     r            ������������������������T     
    long_name    5      Longitude for 2D rectangular grid stored as 1D arrays'        units          degrees_east  �yu�OHDR                                  
   *     �|    �     r            ������������������������R     
    long_name    3      Longitude for 2D irregular grid stored as 1D arrays'        units          degrees_east  J�*OHDR$                                                
   *     �|    �     �            ������������������������S     
    long_name    4      Longitude for 2D rectangular grid stored as 2D array'        units          degrees_east  �U�OHDR$                                                
   *     �|    �     �            ������������������������Q     
    long_name    2      Longitude for 2D irregular grid stored as 2D array'        units          degrees_east  �d�>OHDR    �       �                       
   *     �|   �                 ������������������������+         CLASS          DIMENSION_SCALE "        NAME          lon_T42 +        _Netcdf4Dimid                ����OHDR�    
       
           ?      @ 4 4�     *         �G   �
     P            ������������������������+         CLASS          DIMENSION_SCALE "        NAME          lon_cal +        _Netcdf4Dimid                &    
    long_name          lon_cal/        units          days since 1964-2-28%    	    calendar          365_day%j��OHDRk                      ?      @ 4 4�     *         �G         r            ������������������������(     
    long_name    	      Longitude,        standard_name    	      longitude!        units          degree\        purpose    ?      1-D longitude coordinate referred to by geodesic grid variables  ��%�OHDR�                      ?      @ 4 4�     *         �G    y     r            ������������������������(     
    long_name    	      Longitude,        standard_name    	      longitude!        units          degrees        purpose    V      1-D longitude coordinate referred to by "non-coordinate" (ncd) geodesic grid variables  ���hOHDR                                  
   *     �|   �                 ������������������������+         CLASS          DIMENSION_SCALE "        NAME          lon_grd +        _Netcdf4Dimid                D    
    long_name    %      Longitude grid (typically interfaces)'        units          degrees_east�
��OHDRt                                  
   *     �|    	     r            ������������������������/     
    long_name          Gaussian weights�        purpose    �      Gaussian weights which sum to two for n = 4. These weights are all have floor of 0.0 so should cause SIGFPE when applied to integer types in weighted average.  |��POHDR                      ?      @ 4 4�     *         �G    g�     r            ������������������������P     
    long_name    1      Longitude (typically midpoints), double precision'        units          degrees_east  ��&�OHDR                                  
   *     �|    ��     r            ������������������������P     
    long_name    1      Longitude (typically midpoints), single precision'        units          degrees_east  � l�OHDR                    
   *     �                    ������������������������#     
    long_name          long    �     �        U                                                                                         �ţ�OCHK@        _FillValue                            Η@{?�K�                 OCHKx        purpose    [      Variable of CDL type=long, which is deprecated for int. Included to test back-compatibility[ѵOHDRk    
       ��������    ?      @ 4 4�     +         �G         s            ������������������������6     
    long_name          Least Significant Digit0        purpose          test --lsd switchesp        original_values    K      0.0,0.1,0.12,0.123,0.1234,0.12345,0.123456,0.1234567,0.12345678,0.123456789   ��08OHDR                                   
   *     �|    �     �            ������������������������+         CLASS          DIMENSION_SCALE !        NAME          lsmlev     �      9                            ����BTLF �        c   �        z   �        �   �        �  " �        �   �        �   �           �        $   �        B   �        \   �        v   �        �   �        �   �        �   �        �   �        �  + �        (  + �        S  & �        y   �        �   �        �  & �        �  & �        �  " �          - �        ?  & �        e  & �        �  * �        �  . �          * �        ?  & �        e  1 �        �  0 �        �  * ,�X       OCHK               >        purpose    !      Homebrew level coordinate for LSM)    
    long_name    
      Soil depth         units          meter��OHDR$                                                
   *     �|    t     �            ������������������������E     
    long_name    &      Purpose is to mask a variable like ORO#        units          fraction  �?�OHDR                   *       T                 ������������������������+     
    long_name          the letter a9        purpose          String with known MD5 digestH        MD5_known_checksum           0cc175b9c0f1b6a831c399e269772661/'��OHDR0                              *        	     r            ������������������������.     
    long_name          the letters abc9        purpose          String with known MD5 digestH        MD5_known_checksum           900150983cd24fb0d6963f7d28e17f72  �	OHDR                                  
   *     �|    �	     r            ������������������������J     
    long_name    +      partial mask, partial missing value example@        _FillValue                            Η@{  ���OHDR                                  
   *     �|    c
     r            ������������������������<     
    long_name          partial missing value example@        _FillValue                            Η@{  `�jOHDR                                  
   *     �|    �     r            ������������������������9     
    long_name          all missing values example@        _FillValue                            Η@{  .NOHDR                                  
   *     �|    [     r            ������������������������C     
    long_name    $      offset partial missing value example@        _FillValue                             �y�  ݕ'!OHDR                        
   *     �|   �                 ������������������������3     
    long_name          scalar missing value@        _FillValue                            Η@{                  �Ձ�OHDR�                                  
   *     �|   �                
 �     '�     d�      
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             =$%OHDR1                       
   *     �|   �                 ������������������������M     
    long_name    .      Intended for scalar representation of IEEE NaNb        note    H      20120308 Apparently netCDF ncgen chokes on variable names of nan and NaNk        note2    P      20120330 netCDF ncgen on AIX/bluefire chokes on variable/attribute values of nany        note3    ^      20120625 netCDF ncgen on netCDF 4.1.1 on apparently chokes on variable/attribute values of nan�        note6    �      It is too troublesome to distribute in.cdl with references to NaNs because users always build with old netCDF versions that do not support it. So just comment out nan's for now.@        _FillValue                              �?��D�OHDR                    
   *     �   �                 ������������������������V     
    long_name    7      base date as 6- or 8-digit integer (YYMMDD or YYYYMMDD) 8                                                            ���"BTLF ��  E   �z;! ,   81�! �$   �Q�! 3	   g~"    `�" �  # �Z�" �   f�# �   9�& @   ��' �   BxH' �$  ! �	(    ��( �   ��( �   �~L( �   ���*    Ns_+ G    Z�t+ ?  . ��<, $   ���, �  * �a�, �   ��]- �    <�|- �   7�- 3   ��.    �h�. �  & q<Q/ �   ]��/    j6�0 l   ��2 �   �Qg3 �
   _C�3 u   ���4 _   \��5 Z   7�d6 �   �: �#   �=�: �  $ �{; �   �P�; o"   ��	< �   �w4< r  . *=[< �  . `�W= $  $ �Ҿ� �	   �)� W   ���       OHDR                        
   *     �|   �                 ������������������������+     
    long_name          negative one [                                                                                               @%��OHDR                        
   *     �|   �                 ������������������������H     
    long_name    )      Variable name with pound symbol (invalid) >                                                                  Ty��OHDR                        
   *     �|   �                 ������������������������A     
    long_name    "      Variable name with space (invalid) E                                                                         ԡ~{OHDR                                   
   *     �|   �                 ������������������������/     
    long_name          no missing value    _     Z       +        _Netcdf4Dimid                      h��2OHDR                              *        �     r            ������������������������q     
    long_name    R      Variable contains a one-dimensional array of characters that is not NUL-terminated         units          [chr]  ��$NOHDR$                                            *        �     �            ������������������������r     
    long_name    S      Variable contains a two-dimensional array of characters that are not NUL-terminated         units          [chr]  e��&OHDR�                                *   �    n     r            ������������������������I     
    long_name    *      regular variable, float, packed into short[        purpose    >      Demonstrate that non-rec dim packed vars are handled correctlyB        scale_factor                            ���=@        add_offset                              �B  ��_OHDR     
       ��������            
   +     �   �     
           ������������������������L         DIMENSION_LIST                              D�     �   +        _Netcdf4Dimid                      w�D�OHDR                        
   *     �|   �                 ������������������������"     
    long_name          one d                                                                                                        �ףOHDR                               
   *     �   �                 ������������������������L         DIMENSION_LIST                              D�     �   +        _Netcdf4Dimid                      M7��OHDR                               
   *     �   �                 ������������������������L         DIMENSION_LIST                              D�     �   +        _Netcdf4Dimid                      `u��OHDR     
       ��������            
   +     �   �     
           ������������������������>     
    long_name          one dimensional record variable!        units          kelvin    r�     �              ��Q�OHDRf    
       ��������                
   +     �|    h     s            �������������������������     
    long_name    |      One dimensional record variable with missing data indicated by _FillValue attribute only. No missing_value attribute exists.@        _FillValue                            Η@{   ���OHDR     
       ��������                
   +     �|    v�     s            ������������������������P     
    long_name    1      one dimensional record variable, double precision!        units          second      �I0OHDR     
       ��������                
   +     �|    ZL     R            ������������������������P     
    long_name    1      one dimensional record variable, single precision    ��     Z                              z�OHDR+    
       ��������                
   +     �|    C�     s            ������������������������`     
    long_name    A      one dimensional record variable, single precision, missing values@        _FillValue                            Η@{   -��OHDR{    
       ��������                
   +     �|    �     s            ������������������������h     
    long_name    I      one dimensional record variable, single precision, missing values, scaledB        scale_factor                              �?@        _FillValue                            Η@{   0���OHDR     
       ��������                
   +     �|    3     s            ������������������������X     
    long_name    9      one dimensional record variable, single precision, scaled    ��      P        
              '�=�OCHK    �"     s       @        _FillValue                            Η@{   �(�� OHDR     
       ��������            
   +     �   Y     
           ������������������������M     
    long_name    .      one dimensional record variable to test median    �     Z           �M     9                ��+/OHDR    
       ��������            
   +     �    �     s            ������������������������]     
    long_name    >      one dimensional record variable to test median with _FillValue8        _FillValue                        ���   S�<OHDRi    
       ��������                
   +     �|    o     s            �������������������������     
    long_name    |      One dimensional record variable with missing data indicated by missing_value attribute only. No _FillValue attribute exists.C        missing_value                            Η@{   �XI�OHDR     
       ��������                
   +     �|    �     s            ������������������������U     
    long_name    6      One dimensional record variable with all missing data.@        _FillValue                            Η@{   �d�(OHDR     
       ��������                
   +     �|    �N     R            ������������������������    5E     �      @        _FillValue                              �?    U     Z                        �m�BTLF �          & �        D  + �        o  6 �        �   �        �   �        �   �        �   �        �   �           �        %   �        :   �        T   �        r  . �        �  2 �        �  . �           . �        .  2 �        `  .         �  "        �          �  *          *        ?  .        m  6        �  6        �  *          " 	       %  * 
       O  *        y  *        �  0        �          �   Y�_       OCHK�    
    long_name    �     One dimensional record variable with missing data indicated by a _FillValue attribute that is an array. This can be tested with ncrcat. 20120905: ncgen chokes on _FillValue arrays and produces this error: _FillValue: must be a single (possibly compound) value. Deprecate the array for normal use since it prevents ncgen from completing. Uncommment following line when testing for compatibility with software changes.��Y�OHDRy    
       ��������            +        8     s            ������������������������H     
    long_name    )      one dimensional record variable of string�        NB    �      20131222: HDF4 ncgen fails on this variable: /usr/bin/hncgen -b -o ~/in.hdf ~/nco/data/in.cdl produces error message that "string won't fit in this variable"   ��N�OHDR     
       ��������            
   +     �   8�     
           ������������������������H     
    long_name    )      one dimensional record variable, unsorted         Z           uO     9        	             A�	�OHDRp    
       ��������                
   +     �|    o     s            �������������������������     
    long_name    �      Unsorted, one dimensional record variable with missing data indicated by _FillValue attribute only. No missing_value attribute exists.@        _FillValue                            Η@{   :�g�OHDR                                   
   *     �|   �                 ������������������������L         DIMENSION_LIST                              D�     �        P     9                                U�OHDR�                     *   �   �                 ������������������������G     
    long_name    (      Scalar variable, double, packed as short?       note    %     Original packed value was 1s with scale_factor = 2.0d and add_offset = 1.0d. Unpacked value (netCDF convention) should be 3.0 = 2.0d*1s + 1.0d. Unpacked value (HDF convention) should be 0.0 = 2.0d*(1s-1.0d). NCO algorithms would pack this variable as scale_factor = 0.0d and add_offset = 3.0d.F        scale_factor  ?      @ 4 4�                       @D        add_offset  ?      @ 4 4�                      �?��EOHDR�                     *   �   �                 ������������������������G     
    long_name    (      Scalar variable, double, packed as short?       note    %     Original packed value was 1s with scale_factor = 2.0d and add_offset = 1.0d. Unpacked value (netCDF convention) should be 3.0 = 2.0d*1s + 1.0d. Unpacked value (HDF convention) should be 0.0 = 2.0d*(1s-1.0d). NCO algorithms would pack this variable as scale_factor = 0.0d and add_offset = 3.0d.F        scale_factor  ?      @ 4 4�                       @D        add_offset  ?      @ 4 4�                      �?�G�OHDR�                     *   �                     ������������������������G     
    long_name    (      Scalar variable, double, packed as short?       note    %     Original packed value was 2s with scale_factor = 2.0d and add_offset = 1.0d. Unpacked value (netCDF convention) should be 5.0 = 2.0d*2s + 1.0d. Unpacked value (HDF convention) should be 2.0 = 2.0d*(2s-1.0d). NCO algorithms would pack this variable as scale_factor = 0.0d and add_offset = 5.0d.F        scale_factor  ?      @ 4 4�                       @D        add_offset  ?      @ 4 4�                      �?�rOHDR�                     *   �                    ������������������������G     
    long_name    (      Scalar variable, double, packed as short@       note    &     Original packed value was 1s with scale_factor = 4.0d and add_offset = 3.0d. Unpacked value (netCDF convention) should be 7.0 = 4.0d*1s + 3.0d. Unpacked value (HDF convention) should be -8.0 = 4.0d*(1s-3.0d). NCO algorithms would pack this variable as scale_factor = 0.0d and add_offset = 7.0d.F        scale_factor  ?      @ 4 4�                      @D        add_offset  ?      @ 4 4�                      @G%�POHDR�                                *   �    ��     r            ������������������������F     
    long_name    '      Array variable, double, packed as short]        note    C      Packed value is -32767s, 0s, 1s, 32767s, unpacked is same in doubleF        scale_factor  ?      @ 4 4�                      �?D        add_offset  ?      @ 4 4�                          ��{�OHDR            ?      @ 4 4�     *         �G                    ������������������������!     
    long_name          Pi#        units          fraction 8                                                            MJ��OHDR4    
                     ��������                  �     �       
   +     �|   ��     
                 ������������������������/     
    long_name          Surface pressure!        units          pascal    ;M��OHDR     
       ��������    ?      @ 4 4�     +         �G   ئ     
           ������������������������6     
    long_name          record variable, double    �     Z           �P     9                           ��_�OHDRM    
       ��������              +   �    	     s            ������������������������c     
    long_name    D      record variable, double, packed as short, with double missing valuesJ        purpose    -      Packed version of rec_var_dbl_mss_val_dbl_upk6        _FillValue                       �G        missing_value  ?      @ 4 4�                     8��F        scale_factor  ?      @ 4 4�                   �D        add_offset  ?      @ 4 4�                      @   �h� OHDR�    
       ��������            
   +     �    |     s            ������������������������a     
    long_name    B      record variable, double packed as long, with double missing values�        purpose    e      although not usual, packing doubles into longs (rather than shorts) offers considerable space savings8        _FillValue                        ���G        missing_value  ?      @ 4 4�                     8��F        scale_factor  ?      @ 4 4�                   �D        add_offset  ?      @ 4 4�                      @   �rrOHDR�    
       ��������    ?      @ 4 4�     +         �G    �     s            ������������������������R     
    long_name    3      record variable, double, with double missing values3       purpose         This variable is used to generate the packed variable rec_var_dbl_mss_val_dbl_pck, so its _FillValue should not be out of range, i.e., it should be representable by a short. However, the _FillValue should itself be the same type as the unpacked variable, NC_DOUBLE in this case.D        _FillValue  ?      @ 4 4�                     8��G        missing_value  ?      @ 4 4�                     8��   qr��OHDR>    
       ��������              +   �    �     s            ������������������������b     
    long_name    C      record variable, double, packed as short, with short missing valuesJ        purpose    -      Packed version of rec_var_dbl_mss_val_sht_upk6        _FillValue                       �9        missing_value                       �F        scale_factor  ?      @ 4 4�                   �D        add_offset  ?      @ 4 4�                      @   �w5OHDR�    
       ��������              +   �         s            ������������������������a     
    long_name    B      record variable, double packed as short, with short missing values6        _FillValue                       �F        scale_factor  ?      @ 4 4�                   �D        add_offset  ?      @ 4 4�                      @   ����OHDR�    
       ��������    ?      @ 4 4�     +         �G    �     s            ������������������������R     
    long_name    3      record variable, double, with double missing values3       purpose         This variable is used to generate the packed variable rec_var_dbl_mss_val_sht_pck, so its _FillValue should not be out of range, i.e., it should be representable by a short. However, the _FillValue should itself be the same type as the unpacked variable, NC_DOUBLE in this case.D        _FillValue  ?      @ 4 4�                     8��9        missing_value                       �   ����OHDR�    
       ��������              +   �         s            ������������������������I     
    long_name    *      record variable, double, packed into shortd        purpose    G      Demonstrate that rounding of means of packed data are handled correctlyF        scale_factor  ?      @ 4 4�                �������?D        add_offset  ?      @ 4 4�                      Y@   �|�OHDR     
       ��������                
   +     �|   X�     
           ������������������������5     
    long_name          record variable, float    b     Z           TS     9                                .�&OHDR�    
       ��������                
   +     �|    w     s            ������������������������Q     
    long_name    2      record variable, float, with double missing values@        _FillValue                            Η@{C        missing_value                            Η@{n        note    T      The correct average of this variable is 5.0. The correct sum of this variable is 35.   緳�OHDR     
       ��������                
   +     �|    #%     s            ������������������������P     
    long_name    1      record variable, float, with float missing values    T     N           �S     9         )hl�FSSE �        �     �   �   �   �	   �     �   
  �     �     �     �   � %   ���)OHDR-    
       ��������                
   +     �|     "     s            ������������������������b     
    long_name    C      record variable, float, with float missing values in every position@        _FillValue                            Η@{   Y}s0OHDR     
       ��������                
   +     �|    �<     g            ������������������������j     
    long_name    K      record variable, float, with float missing values in every position but one                   pe�BTLF �x�� �  * ��� �   ��,� �   ��� �
   ~��� 0   �v�� -"    BUQ� +   ��� �   ^k�� A   ׅ9� J   ~�r� ?  & L�� �   ��� �   H��� �   ��>� �   �\��    ���� %   g8� �   �T�� :   ���� �
   ɤ�� O  ! �O� �!   e�� �   �7:� �   �	|� �  . <@�� �  & q<Q/ �   ]��/    j6�0 l   ��2 �   �Qg3 �
   _C�3 u   ���4 _   \��5 Z   7�d6 �   �: �#   �=�: �  $ �{; �   �P�; o"   ��	< �   �w4< r  . *=[< �  . `�W= $  $ �Ҿ� �	   �)� W   ���       OHDR5    
       ��������                
   +     �|    #     s            ������������������������j     
    long_name    K      record variable, float, with float missing values in every position but two@        _FillValue                            Η@{   �ArzOHDR^    
       ��������                
   +     �|    y#     s            ������������������������R     
    long_name    3      record variable, float, with integer missing values@        _FillValue                             �y�;        missing_value                        ���   �L��OHDR�    
       ��������              +   �    �#     s            ������������������������H     
    long_name    )      record variable, float, packed into shortd        purpose    G      Demonstrate that rounding of means of packed data are handled correctlyB        scale_factor                            ���=@        add_offset                              �B   3{:OHDR[    
       ��������            
   +     �    _$     s            ������������������������S     
    long_name    4      record variable, integer, with double missing values8        _FillValue                        ���G        missing_value  ?      @ 4 4�                     8��   y��DOHDRV    
       ��������            
   +     �    	)     s            ������������������������R     
    long_name    3      record variable, integer, with float missing values8        _FillValue                        ���C        missing_value                             �y�   ߱z:OHDR    
       ��������            
   +     �    �%     s            ������������������������T     
    long_name    5      record variable, integer, with integer missing values8        _FillValue                        ���   V��OHDR�    
       ��������              +   �    	&     s            ������������������������B     
    long_name    #      Array packed with scale factor only�        note    �      Original packed value was 1s..10s with scale_factor = 10.0d no add_offset. Unpacked value should be 10.0 = 10.0d*1s + 0.0d through 100 = 10.0d*1s + 0.0d. Average value should be 55.F        scale_factor  ?      @ 4 4�                      $@   ���OHDRT                                  
   *     �|    �&     �            ������������������������+         CLASS          DIMENSION_SCALE         NAME          rlev +        _Netcdf4Dimid                I        purpose    ,      Monotonically decreasing coordinate pressure  8�fOHDR*                                  
   *     �|    |&     r            ������������������������%     
    long_name          Height         units          meterU        purpose    8      Height stored with a monotonically decreasing coordinate  Â3OHDR                        
   *     �|   ,                 ������������������������.     
    long_name          scalar variable#        units          fraction /                                                   ?���BTLF                  :          V          k          �          �  $        �           �  $           $        $  $        H  $        l          �          �          �          �               !       .    "       G    #       `    $       y    %       �    &       �    '       �    (       �    )       �   " *       !  & +       :!   ,       X!   -       m!   .       �!   �TU�     �          �   Y�_       OHDR�                     *   �   0                 ������������������������>     
    long_name          scalar variable, double, packedQ        purpose    4      Packed version of number with ncdiff subtraction bugF        scale_factor  ?      @ 4 4�                   �D        add_offset  ?      @ 4 4�                      @TբEOHDR                      *   �   2                 ������������������������$     
    long_name          short l                                                                                                                ��:OHDR$    
              ��������           �'     �       
   +     �|   �J     
              �������������������������     
    long_name    e      two dimensional record variable stored in td (time,dgn) order (dgn means degenerate, i.e., of size 1)    �[��OHDRP4    
                     ��������                          
   +     �    �=     �                      ������������������������@     
    long_name    !      three dimensional record variable'        units          watt meter-28        _FillValue                        �������OHDR                        
   *     �|   4                 ������������������������$     
    long_name          three b                                                                                                      E(UOHDR4    
                     ��������                  k�     �       
   +     �|   a     
                 ������������������������@     
    long_name    !      three dimensional record variable'        units          watt meter-2    <��OHDRL4                                                              
   *     �|          �            ������������������������     
    long_name    `      three dimensional variable with CCM coordinate convention C=[lat,lev,lon], Fortran=(lon,lev,lat)#        units          fraction  ?h�qOHDRO4                                                              
   *     �|    �     �            �������������������������     
    long_name    c      three dimensional variable with COORDS coordinate convention C=[lev,lat,lon], Fortran=(lon,lat,lev)#        units          fraction  �ʜgOHDRw4    
                     ��������                  $     �          +         �G   Pm     
                 ������������������������O     
    long_name    0      three dimensional record variable of type double'        units          watt meter-2D        _FillValue  ?      @ 4 4�                     �X�    �_EOHDR\4    
                     ��������                          
   +     �    �     �                      ������������������������L     
    long_name    -      three dimensional record variable of type int'        units          watt meter-28        _FillValue                        ����(qH�OHDRL4    
                     ��������                            +   �    �      �                      ������������������������@     
    long_name    !      three dimensional record variable'        units          watt meter-26        _FillValue                       ����vLOHDR�    
       ��������    ?      @ 4 4�     +         �G  L �W     �          N ������������������������+         CLASS          DIMENSION_SCALE         NAME          time +        _Netcdf4Dimid                #    
    long_name          time?        units    $      days since 1964-03-12 12:09:00 -9:00'    	    calendar    	      gregorian%        bounds    	      time_bnds   �]�OHDR $    
              ��������           �Y     S       
   +     �|   @�     
              ������������������������@         purpose    #      Cell boundaries for time coordinate     !     j                           Pm�OHDR $    
              ��������           GZ     S       
   +     �|   x�     
              ������������������������F     
    long_name    '      Record variable of longitude coordinate    �!     j        	             �� OHDR�                      ?      @ 4 4�     *         �G   �                 ������������������������+         CLASS          DIMENSION_SCALE '        NAME          time_udunits +        _Netcdf4Dimid                ;        units           hours since 1900-01-01 00:00:0.01        delta_t          0000-00-00 06:00:0.0Q        purpose    4      The dates specified in this variable are ~1999-12-08L��OHDR            ?      @ 4 4�     *         �G                    ������������������������0         units          days since 2013-01-01%    	    calendar          360_day '                                           a�
�OHDR            ?      @ 4 4�     *         �G                    ������������������������0         units          days since 2013-01-01%    	    calendar          365_day '                                           7��[OCHKL        DIMENSION_LIST                              D�        ~1��FSSE �      �  ;    "� OHDR            ?      @ 4 4�     *         �G                     ������������������������0         units          days since 2013-01-01%    	    calendar          366_day '                                           � C�OHDR            ?      @ 4 4�     *         �G   (                 ������������������������0         units          days since 2013-01-01'    	    calendar    	      gregorian %                                         猅�OHDR            ?      @ 4 4�     *         �G   0                 ������������������������0         units          days since 2013-01-01$    	    calendar          julian (                                            B
+�BTLF 9��b H  $ �bc �   e��c �   �|�c �  " ���e �   CH^f t   %�uf �   8k�g 
   k��h 3   i(�h �   A/?i $   ��i V   o��i �   ��i Y$   �KWj m
   �sNk �"  " ��ll W
   ��l �	   D�l �   @�0m �   �n V   On    �mVn X!   {Fo �	   s&o �   �Ho S  & �y�o �    d�;p   " �8�p ,   T@-q �   V��q T   �`2r �   �7r �
   �l�r    $ ��s `  . Z$�s �   ́lt p   ��t _   ��v m   %��v O  * ��Iw �   ��Yx �"   �	�z �   j� �	   �)� W   ���       OHDR            ?      @ 4 4�     *         �G   8                 ������������������������0         units          days since 2013-01-01 R                                                                                      ��;�OHDR+    
       ��������                
   +     �|    ,     s            ������������������������*     
    long_name          Temperature!        units          kelvinO        hieght    3      Leave hieght mispelled for NCO User's guide example   z���OHDR    
       ��������    ?      @ 4 4�     +         �G    dB     s            ������������������������T     
    long_name    5      Temperature stored as double precision floating point!        units          kelvin   k�SOHDR     
       ��������                
   +     �|    �,     s            ������������������������T     
    long_name    5      Temperature stored as single precision floating point!        units          kelvin   H�OHDR                        
   *     �|   @                 ������������������������"     
    long_name          two d                                                                                                        e��OHDR$    
              ��������           �,     �       
   +     �|   @�     
              ������������������������>     
    long_name          two dimensional record variable'        units          watt meter-2    i�W�OHDR $    
              ��������                   +       x�     
              ������������������������H     
    long_name    )      two dimensional record variable of string    1>     j           �[     9         ���OHDR $                                                
   *     �|    �>     �            ������������������������7     
    long_name          two dimensional variable#        units          fraction             ��dOOHDR $    
              ��������           ?     �       
   +     �|   ��     
              ������������������������\     
    long_name    =      two dimensional record variable stored in tx (time,lon) order 	             a���OHDR(D    
                            ��������                         |)     �       
   +     �|   ��     
                    ������������������������g     
    long_name    H      four dimensional record variable stored in txyz (time,lon,lat,lev) order    x$OHDR $    
              ��������            *     �       
   +     �|   0�     
              ������������������������\     
    long_name    =      two dimensional record variable stored in ty (time,lat) order 	             ��q�OHDR $    
              ��������           �*     �       
   +     �|   h�     
              ������������������������\     
    long_name    =      two dimensional record variable stored in tz (time,lev) order 	              J�BOHDR     
       ��������                
   +     �|    �]     R            ������������������������/     
    long_name          Zonal wind speed)        units          meter second-1    �     Z                ���9OHDR            ?      @ 4 4�     *         �G   \                 ������������������������7     
    long_name          Unpacked scalar variable    �            5                                                         ���6BTLF 0       �   1       �!   2       �!   3       �!   4       �!    5       "   6       -"    7       M"  " 8       o"   9       �"   :       �"  " ;       �"  " <       �"   =       #   >       )#   ?       F#   @       c#   A       }#   B       �#   C       �#   D       �#   E       �#   F       $   G       $   H       ,$   I       C$   J       Y$   K       t$  ! L       �$  ! M       �$   N       �$   O       �$  ! ^�¹     �   Y�_       OCHK       note    �      Unpacked value is 3.0d0, upk=unpack(pck)= 2.0d0*1s + 1.0d0 = 3.0d0. Packing this variable should create an NC_SHORT scalar = 0s with packing attribute add_offset=3.0d and either no scale_factor (ncap) or scale_factor = 0.0d (ncpdq).|A6OHDR�                      ?      @ 4 4�     *         �G    (+     r            ������������������������-     
    long_name          Unpacked array�        note    �      Unpacked value is -32767.d, 0.d, 1.d, 32767.d, packed is same in short. Packing algorithm should yield an NC_SHORT array = [] with packing attributes scale_factor=1.0d, add_offset=0.0d  �Eu?OHDR     
       ��������                
   +     �|    \^     R            ������������������������4     
    long_name          Meridional wind speed)        units          meter second-1    �(     Z            q�%�OHDR(                       
   *     �|   �                 ������������������������k     
    long_name    L      Floating point number with exponent ending in zero to test sng_trm_trl_zro()C        att_eminusten                            ��.���POHDR                        
   *     �|   �                 ������������������������4     
    long_name          Scalar with value 0.5@        _FillValue                            Η@{                 �n�OHDR                                   
   *     �|    �+     r            ������������������������&     
    long_name          0.5,0.5@        _FillValue                            Η@{                 f>�cOHDR                                 *   �    �^     Q            ������������������������+     
    long_name          17000, 170006        _FillValue                       ��    �E     Z                 �l�OHDR                    
   *     �   �                 ������������������������8     
    long_name          scalar integer equal to 18        _FillValue                        ����                             �]��OHDR                                  
   *     �|    �H     r            ������������������������C     
    long_name    $      one regular value, one missing value@        _FillValue                            Η@{  �|�]OHDR                               
   *     �    �_     Q            ������������������������)     
    long_name    
      1, mss_val8        _FillValue                        ����    I     Z               �%�OHDR                               
   *     �    �_     Q            ������������������������#     
    long_name          1, 18        _FillValue                        ����    qI     Z        	             �4]�OHDR                                   
   *     �|    C`     Q            ������������������������S     
    long_name    4      Variable for 2D rectangular grid stored as 1D arrays    �B     Z                           �4�OHDR                                   
   *     �|    �`     Q            ������������������������Q     
    long_name    2      Variable for 2D irregular grid stored as 1D arrays    1C     Z                             Rr&FOHDR $                                                
   *     �|    �`     Q            ������������������������R     
    long_name    3      Variable for 2D rectangular grid stored as 2D array    �C     j             "hs�OHDR $                                                
   *     �|    6a     Q            ������������������������P     
    long_name    1      Variable for 2D irregular grid stored as 2D array    �C     j              ?x�OHDR$                                                
   *     �|    _D     �            ������������������������G     
    long_name    (      Float field for testing masks and wheres#        units          fraction  �̑�OHDR                       
   *     �|   T                 ������������������������S     
    long_name    4      Variable and attribute names include dash charactersA        att_nm-dash                            Η@{�{��OHDR    
       ��������                
   +     �|    �D     �            ������������������������*     
    long_name          Temperature�        purpose    v      Array containing _FillValue at some locations, out-of-range values at other locations, and valid data in the remainder@        _FillValue                             �y�?    
    valid_min                              4C?    
    valid_max                              �C   M5�vOHDR                                   
   *     �|    �a     Q            ������������������������.     
    long_name          Gaussian weight#        units          fraction    �E     Z                       +��$OHDR                                   
   *     �|   `                 ������������������������1     
    long_name          all values are one    =F     Z       +        _Netcdf4Dimid                    ��OHDRK4    
                     ��������                  �F     �       
   +     �|   0!     
                 ������������������������)     
    long_name    
      wind speed)        units          meter second-1@        _FillValue                             �y�    ����OHDRY                                  
   *     �|   p-                 ������������������������+         CLASS          DIMENSION_SCALE         NAME          wvl +        _Netcdf4Dimid                )    
    long_name    
      Wavelength         units          meterE�2OHDR*                                  
   *     �|    +G     r            ������������������������%     
    long_name          Height         units          meterU        purpose    8      Height stored with a monotonically increasing coordinate  �o�OHDR                        
   *     �|   �-                 ������������������������#     
    long_name          zero c                                                                                                       ��EGOHDR8                     !               
   �     �            ������������������������+         CLASS          DIMENSION_SCALE Z        NAME    @      This is a netCDF dimension but not a netCDF variable.         2 +        _Netcdf4Dimid                  ¼�=OHDR8                     !               
    F�     �            ������������������������+         CLASS          DIMENSION_SCALE Z        NAME    @      This is a netCDF dimension but not a netCDF variable.         5 +        _Netcdf4Dimid                  ��IOHDR8                     !               
    C�     �            ������������������������+         CLASS          DIMENSION_SCALE Z        NAME    @      This is a netCDF dimension but not a netCDF variable.        26 +        _Netcdf4Dimid             	     ��%�OHDR8    P       P          !               
   _�     �            ������������������������+         CLASS          DIMENSION_SCALE Z        NAME    @      This is a netCDF dimension but not a netCDF variable.        80 +        _Netcdf4Dimid                  fBOHDR8                     !               
   ��     �            ������������������������+         CLASS          DIMENSION_SCALE Z        NAME    @      This is a netCDF dimension but not a netCDF variable.         8 +        _Netcdf4Dimid                  8r��OHDR8                     !               
   �     �            ������������������������+         CLASS          DIMENSION_SCALE Z        NAME    @      This is a netCDF dimension but not a netCDF variable.         2 +        _Netcdf4Dimid                  +���OHDR8                     !               
   �     �            ������������������������+         CLASS          DIMENSION_SCALE Z        NAME    @      This is a netCDF dimension but not a netCDF variable.         4 +        _Netcdf4Dimid                  s�tZOCHK    �$     Q       \        DIMENSION_LIST                              D�           D�          N��GCOL                        �                    �                    �                    
�                    
�                    ��                    s�                   s�     	              
�      
              s�                   
�                    ��                    s�                   
�                    
�                    
�                    s�                   t�                    t�                    ��                   
�                    
�                    ��                    
�                    
�                    t�                    
�                    t�                    ��                    s�                   s�                    
�      !              s�     "              
�      #              ��      $              
�      %              
�      &              ��      '              ��      (              s�     )              s�     *              s�     +              s�     ,              *�     -              s�     .              s�     /              n�     0              �      1              ��     2              &�      3              &�      4              ��     5              s�     6              s�     7              ��     8              ��      9              ��      :              s�     ;              s�     <              
�      =              s�     >              
�      ?              t�      @              s�     A              
�      B              t�      C              ��      D              s�     E              s�     F              ��      G              ��      H              ��     I              
�      J              �      K              t�      L              t�      M              t�      N              t�      O              :�     P              g�      Q              g�      R              
�      S              
�      T              ��      U              
�      V              
�      W              ��      X              
�      Y              
�      Z              :�     [              
�      \              ��      ]              ��     ^              
�      _              
�      `              t�      a              t�      b              t�      c              g�      d              g�      e              
�      f              
�      g              ��      h              
�      i              
�      j              ��      k              ��      l              ��     m              ��      n              ��      o              ��      p              s�     q              
�      r              
�      s              ��      t              t�      u              ��      v              ��      w              ��      x              ��      y              
�      z              ��      {              ~�     |              &�      }              &�      ~              ~�                   ��      �              s�     �              
�      �              
�      �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              ��     �              ��      �              s�     �              s�     �              
�      �              s�     �              
�      �              ��      �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     �              s�     OCHK   ��            l     0   REFERENCE_LIST 6     dataset        dimension                        �              ��OCHK   @�             l     0   REFERENCE_LIST 6     dataset        dimension                        �             ��ݰOCHK    �     Q       \        DIMENSION_LIST                              D�           D�          �d�OCHKl         DIMENSION_LIST                              D�           D�           D�        �3�gBTHD 	      d(�     
 
       ���  OCHKL        DIMENSION_LIST                              D�        �;i�FSSE K�     
  �    s �    ٻ��   OCHK    2H     S       l        DIMENSION_LIST                              D�     
      D�           D�            h���FRHP               ���������      W                           	                                                      (  �}       2���BTHD 	      d(p;     	 	       � 1�          OCHKL        DIMENSION_LIST                              D�        V�
�OCHK\        DIMENSION_LIST                              D�     %      D�     &   �9�OOCHKL        DIMENSION_LIST                              D�     J   MHЏOCHK   |�            l     0   REFERENCE_LIST 6     dataset        dimension                        x�              ���FHIB �          �\     P     ������������������-�OCHK   ��             +        _Netcdf4Dimid                ����                 D�           D�        �O5�OCHK    9P     Q       L        DIMENSION_LIST                              D�     �     ����                                OCHK                |        DIMENSION_LIST                              D�     @      D�     A      D�     B      D�     C   +        _Netcdf4Dimid                sI3E                             OCHKl         DIMENSION_LIST                              D�     !      D�     "      D�     #   ^	�kOCHK   ��     
      L        DIMENSION_LIST                              D�     )   +        _Netcdf4Dimid                ��~9                               OCHK    J�     Q       L        DIMENSION_LIST                              D�     '     w�4OCHK    W@     Q       L        DIMENSION_LIST                              D�     G     ����                                OCHK    UW     R       L        DIMENSION_LIST                              D�     (      �u#OCHKL        DIMENSION_LIST                              D�     +   w^��OCHKL        DIMENSION_LIST                              D�     ,   |��LBTHD       d(p9     	 	       ,L=         OCHKL        DIMENSION_LIST                              D�     *   �H?LOCHK    ��������h       l     0   REFERENCE_LIST 6     dataset        dimension                        ��             j�#@OCHKL        DIMENSION_LIST                              D�     0   쿝n                       OCHK    ��������       l     0   REFERENCE_LIST 6     dataset        dimension                        �              5��OCHK    >     V             \        DIMENSION_LIST                              D�     .      D�     /   ��wOCHK    ��������@      �     0   REFERENCE_LIST 6     dataset        dimension                        ��              ��             ��             ����OCHKL        DIMENSION_LIST                              D�     I   �!�
OCHK    �W     S       l        DIMENSION_LIST                              �-           �-           �-            �*�     OCHKL        DIMENSION_LIST                              D�     1   *{ 4OCHK    ?     V             \        DIMENSION_LIST                              D�     6      D�     7   ��/           OCHK    �>     Q       \        DIMENSION_LIST                              D�     3      D�     4     ���mOCHKL        DIMENSION_LIST                              D�     �   +        _Netcdf4Dimid                ٓ��       OCHK    b?     Q       L        DIMENSION_LIST                              D�     8     thaOCHK    L     R       L        DIMENSION_LIST                              D�     �      `�"nOCHKL        DIMENSION_LIST                              D�     �   *�OCHK    �L     R       L        DIMENSION_LIST                              D�     �      f��                   OCHK    �?     Q       L        DIMENSION_LIST                              D�     9     ���;OCHK     C     Q       \        DIMENSION_LIST                              D�     V      D�     W     ���OCHK\        DIMENSION_LIST                              D�     Y      D�     Z   S��BTHD       d(�     
 
       LX6�OCHK    @     S       \        DIMENSION_LIST                              D�     E      D�     F       ��X9OCHK    ��������        �     0   REFERENCE_LIST 6     dataset        dimension                        ��              Q�              �             \LW OCHK    �@     Q       L        DIMENSION_LIST                              D�     H     ���OCHK    �E     Q       L        DIMENSION_LIST                              D�     c     ��HvOCHK    �G     Q       L        DIMENSION_LIST                              D�     n     ����OCHK    :H     Q       L        DIMENSION_LIST                              D�     o      �D�FSHD  }                             P x (        ��     %       %       ���FSSE �V     � l    �1	� OCHKL        DIMENSION_LIST                              D�     K   �F�OCHKL        DIMENSION_LIST                              D�     L   ��]OCHK\        DIMENSION_LIST                              D�     N      D�     O   ��ÿOCHK    �C     Q       L        DIMENSION_LIST                              D�     \     �T                                OCHK    B     Q       L        DIMENSION_LIST                              D�     P     =���OCHK    �B     Q       \        DIMENSION_LIST                              D�     S      D�     T     �J��                OCHK    ^B     Q       L        DIMENSION_LIST                              D�     Q     ����OCHK    F     Q       L        DIMENSION_LIST                              D�     d     ����OCHK   X�             �     0   REFERENCE_LIST 6     dataset        dimension                        ��              f�             �              ��                           �Zz�                                OCHK    D     Q       L        DIMENSION_LIST                              D�     ]     ���~OCHK    ��������       �     0   REFERENCE_LIST 6     dataset        dimension                        ��             !�             O�            [�w0                              OCHK    �F     Q       \        DIMENSION_LIST                              D�     i      D�     j     y�oOCHK    �F     Q       L        DIMENSION_LIST                              D�     k     t":�OCHK    GG     Q       L        DIMENSION_LIST                              D�     l     �i�DOCHK                �  	   0   REFERENCE_LIST 6     dataset        dimension                        ��              ��              �              �              R�             ^�             �K
            OCHK    TF     Q       \        DIMENSION_LIST                              D�     f      D�     g     =�R�OCHK    rJ     Q       L        DIMENSION_LIST                              D�     x     �T�FRHP               ��������Q      K�                          
                                                      (  �      g�QlOCHKL        DIMENSION_LIST                              D�     z   ��IHOCHK   `�             +        _Netcdf4Dimid                �G�   OCHK    �G     Q       L        DIMENSION_LIST                              D�     m     Z.�VOCHK    .I     Q       L        DIMENSION_LIST                              D�     t     R*�OCHK    I     Q       L        DIMENSION_LIST                              D�     u     ���OCHK    �I     Q       L        DIMENSION_LIST                              D�     v     �
�8BTHD       d(p5     	 	       �[K�      OCHK    �H     R       L        DIMENSION_LIST                              D�     p      ����OCHK    �H     Q       \        DIMENSION_LIST                              D�     r      D�     s     �щPOCHK    �J     Q       L        DIMENSION_LIST                              D�     {     ;F��OCHK    �K     R       L        DIMENSION_LIST                              D�     �      +}W                               OCHK    K     Q       \        DIMENSION_LIST                              D�     }      D�     ~     K�ۨOCHK+        _Netcdf4Dimid                5��   OCHK    !J     Q       L        DIMENSION_LIST                              D�     w     �|?1OCHK   �            |     0   REFERENCE_LIST 6     dataset        dimension                        ��              y-             b��OCHK    ��������       |     0   REFERENCE_LIST 6     dataset        dimension                        a,             y-            �︣OCHK    eK     Q       L        DIMENSION_LIST                              D�          Gۺ.FSSE W     � -    o�˘ BTLF  �   \     қ-     L      L�  /   y     �>q b    b     ��# �   @     �$ �    k     �V�k b   +  	   e>� �   �     ��� �   �     �)m�    L     c����Zڵ                                                                                                                                                                                                                                                                                                                                            BTLF 	     L       b    b      �    k      /   y      �   �      �   \      �   �      �   @         L      b   +  	   �A_u                                                                                                                                                                                                                                                                                                                                                                                    OCHK    �M     R       L        DIMENSION_LIST                              D�     �      �5�OCHK    -N     R       L        DIMENSION_LIST                              D�     �      ���BOCHK    N     R       L        DIMENSION_LIST                              D�     �      ��+mOCHKL        DIMENSION_LIST                              D�     �   #]E�OCHKL        DIMENSION_LIST                              D�     �   {��OCHK    Q     R       L        DIMENSION_LIST                              D�     �      ����OCHK    hQ     R       L        DIMENSION_LIST                              D�     �      N$�OCHK    �Q     R       L        DIMENSION_LIST                              D�     �      blmOCHKL        DIMENSION_LIST                              D�     �   D�*m    OCHK    �L     R       L        DIMENSION_LIST                              D�     �      q!OCHK    PM     R       L        DIMENSION_LIST                              D�     �      ����OCHKL        DIMENSION_LIST                              D�     �   Ϯ:DOCHK    KX     Q       l        DIMENSION_LIST                              �-           �-           �-          ��*OCHK    �X     Q       l        DIMENSION_LIST                              �-           �-           �-          �ˇ�OCHK    �X     S       l        DIMENSION_LIST                              �-     #      �-     $      �-     %       ���OCHKL        DIMENSION_LIST                              �-     W   �T%t   OCHKL        DIMENSION_LIST                              D�     �   E@)OCHK    �O     R       L        DIMENSION_LIST                              D�     �      ��MOCHK    ��������       |     0   REFERENCE_LIST 6     dataset        dimension                        E�             K             �)�(OCHK    �P     S       l        DIMENSION_LIST                              D�     �      D�     �      D�     �       �E��                                OCHK    #O     R       L        DIMENSION_LIST                              D�     �      g�jOCHK    R     R       L        DIMENSION_LIST                              D�     �      ��mOCHK    ^R     R       L        DIMENSION_LIST                              D�     �      8��OCHK    �R     R       L        DIMENSION_LIST                              D�     �      ��OCHK    S     R       L        DIMENSION_LIST                              D�     �      ���OCHK    �S     R       L        DIMENSION_LIST                              D�     �      u��OCHK    @Y     Z                l        DIMENSION_LIST                              �-     )      �-     *      �-     +   ��OCHK    �Y     Z                l        DIMENSION_LIST                              �-     /      �-     0      �-     1   5�)�OCHK\        DIMENSION_LIST                              �-     3      �-     4   ͼ �OCHK\        DIMENSION_LIST                              �-     6      �-     7   ����BTHD 	      d(p7     	 	       ���      OCHK    T     R       L        DIMENSION_LIST                              D�     �      h��[OCHK    jT     R       L        DIMENSION_LIST                              D�     �      �sc;OCHK    �T     R       L        DIMENSION_LIST                              D�     �      �I�MOCHK    U     R       L        DIMENSION_LIST                              D�     �      �O��OCHK    `U     R       L        DIMENSION_LIST                              D�     �      V�y_OCHK    �U     R       L        DIMENSION_LIST                              D�     �      ���(OCHK    �     @       +        _Netcdf4Dimid                 ����OCHK   ��     
      L        DIMENSION_LIST                              D�     �   ��tOCHK    VV     R       L        DIMENSION_LIST                              �-           ��uOCHK    �V     R       L        DIMENSION_LIST                              �-           >�OCHK    �V     Q       L        DIMENSION_LIST                              �-          ��6�OCHK               l     0   REFERENCE_LIST 6     dataset        dimension                        �             =�d�OCHK    KW     S       \        DIMENSION_LIST                              �-           �-            ~�J�OCHK   ��            |     0   REFERENCE_LIST 6     dataset        dimension                        y�              Ɔ            ��DVOCHKL        DIMENSION_LIST                              �-     Y   ^+qj         OCHK    V     R       L        DIMENSION_LIST                              �-           8�G�OCHK    �\     S       |        DIMENSION_LIST                              �-     M      �-     N      �-     O      �-     P       �:��OCHK    ]     S       \        DIMENSION_LIST                              �-     R      �-     S       �3�@OCHK    f]     S       \        DIMENSION_LIST                              �-     U      �-     V       �ՆdOCHK    ^     Q       L        DIMENSION_LIST                              �-     X     ���OCHK    �^     Q       L        DIMENSION_LIST                              �-     Z     !m��  OCHK    �Z     R       L        DIMENSION_LIST                              �-     8      O�oOCHK    >[     R       L        DIMENSION_LIST                              �-     :      ݣ��OCHK    �[     S       \        DIMENSION_LIST                              �-     <      �-     =       �笶                              GCOL                        s�                   s�                   s�                   w~                   s�                   s�                   �                    s�     	              s�     
              
�                    s�                   
�                    ��                    s�                   s�                   
�                    s�                   
�                    ��                    
�                    
�                    t�                    
�                    t�                    ��                    t�                    t�                    
�                    t�                    
�                    ��                     s�     !              s�     "              
�      #              s�     $              
�      %              ��      &              s�     '              s�     (              
�      )              s�     *              
�      +              ��      ,              s�     -              s�     .              
�      /              s�     0              
�      1              ��      2              s�     3              s�     4              :�     5              s�     6              s�     7              ��      8              s�     9              s�     :              s�     ;              s�     <              s�     =              t�      >              s�     ?              s�     @              t�      A              
�      B              
�      C              t�      D              s�     E              s�     F              ��      G              s�     H              s�     I              ��      J              s�     K              ��      L              
�      M              s�     N              ��      O              
�      P              t�      Q              s�     R              s�     S              
�      T              s�     U              s�     V              t�      W              s�     X              ��      Y              s�     Z              
�      [              
�      \              
�      ]              
�      ^              
�      _              g�      `              g�      a              
�      b              
�      c              ��      d              
�      e              
�      f              ��      g              
�      h              
�      i              ��      j              s�     k              
�      l              
�      m              s�     n              s�     o              
�      p              s�     q              
�      r              ��      s              t�              (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              OCHK    �W     Z                l        DIMENSION_LIST                              �-           �-           �-        Pp�OCHK\        DIMENSION_LIST                              �-     ?      �-     @   ���7OCHK    \     Q       \        DIMENSION_LIST                              �-     B      �-     C     �2IOCHK    m\     S       \        DIMENSION_LIST                              �-     E      �-     F       �6��FHDB �         ��oR�       e_dbl��      �       e_flt�      �       fl_dmn&�      �       fl_nm��      �       	fl_nm_arr��      �       	fl_nm_rec��      �       fll_val��      �       fll_val_mss_val��      �       	float_var	�      �       four�      �       four_dmn_rec_var!�      �       gZ�      �       	gds_3dvarf�      �       gds_crd��      �       gds_var�      �       gds_var_ncd��      �       gwl�      �       gw_T42x�                      OCHK   0�            +        _Netcdf4Dimid                �.6�OCHK   8�            +        _Netcdf4Dimid                r�                                 OCHK    �Z     R       L        DIMENSION_LIST                              �-     9      ��T�OCHKL        DIMENSION_LIST                              �-     _   ����OCHKL        DIMENSION_LIST                              �-     `   �<�OCHK\        DIMENSION_LIST                              �-     b      �-     c   a6�OCHK\        DIMENSION_LIST                              �-     e      �-     f   nѕ�OCHK    �a     Q       \        DIMENSION_LIST                              �-     h      �-     i     ��GOCHK         
      L        DIMENSION_LIST                              �-     j   +        _Netcdf4Dimid                ��G�    OCHKL        DIMENSION_LIST                              �-     [   ���OCHKL        DIMENSION_LIST                              �-     k   ����OCHKL        DIMENSION_LIST                              �-     l   ��ӒOCHK    )b     S       l        DIMENSION_LIST                              �-     p      �-     q      �-     r       i��OCHK    |b     Q       L        DIMENSION_LIST                              �-     s     
:��FHIB �          ؆     ؄     ؂     ؀     �~     �|     T     �?     �x     �p     �l     �h     �`     �������������������������cOCHK                +        _Netcdf4Dimid                ﳚ#                                OCHK    P_     Q       L        DIMENSION_LIST                              �-     \     '�`OCHKL        DIMENSION_LIST                              �-     ]   �-nOCHKL        DIMENSION_LIST                              �-     ^   �~�OCHK   �            , 2   0   REFERENCE_LIST 6     dataset        dimension          -       -       D              �             ��              ��              ��              ��              ��              ��             ��              !�             l�              ��              ��              !�              ��              \�              h�              $              D             u             N             x2             �3             MY            �            W�            }�             Ռ            0�            ��            �            ��             ��            ت            ��             	�             !�             :�             F�             j�             v�             ��             ��             ��             ��            Q�sOCHK   d            � ,   0   REFERENCE_LIST 6     dataset        dimension          (       (       D             �             ��             ��             ��             ��             ��              ��              !�             ��             ��             $             D            �	             *             ;             u            �                                       )             U+             �.             |V             MY            �            W�            }�            Ռ            0�            ��            �            [�            ��            ��            �             j�            v�            ��            ��            kp7FHDB �         `�(     DIMENSION_LIST                              D�     y        _Netcdf4Dimid                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   FHDB �         ���       char_var٥      �       char_var_nul�      �       char_var_space�      �       
cnv_CF_crd��      �       
cnv_CF_ncl��      �       cnv_CF_ncl_var_1|�      �       cnv_CF_ncl_var_2�      �       date߱      �       date_int�      �       date_rec��      �       dgn�      �       dgn_vary�      �       
double_var��      �       double_var2��      �       dps_dry��      �       dps_ttl��      �       dps_wet��                FRHP               ���������      �V                           	                                                      (  ��       ��GhFSHD  �                             P x (        ��                   �%FSHD  �                             P x (        �                   ⼆jOCHK   ��     
      +        _Netcdf4Dimid                0�
OCHK+        _Netcdf4Dimid                �w�     OCHK   �     
      � M   0   REFERENCE_LIST 6     dataset        dimension          G       G       �              ��              ��              ��              ��              |�              �              ߱              ��              ��              !�              f�              9             `0             �4             �5             7             8             &9             ]:             �;             X=             d>             �?             �@             )B             G             �H             �I             MY             \Z             h[             �]             T`             c             Ue             g             �i             �k             �l             yn             �o             +q             7t             xu             �v             �x             z             r{             �|             Ɔ             �             W�             0�             ��             �             O�             [�             �             H�             X�             p�             ��             ��             ��             ت             �             �             ��             ��             ��             �&VFHDB �          b�S� 
    long_name    -      Intended for array representation of IEEE NaN     note    H      20120308 Apparently netCDF ncgen chokes on variable names of nan and NaN     note2    P      20120330 netCDF ncgen on AIX/bluefire chokes on variable/attribute values of nan     note3    ^      20120625 netCDF ncgen on netCDF 4.1.1 on apparently chokes on variable/attribute values of nan     note4    �      If your NCO build fails because your version of netCDF does not support nan, then cd to the directory that contains the file nco/data/in.cdl and run the command in note5 first and then try to build again     note5    A      sed -e 's/nan;/1.0f;/' in.cdl > foo.cdl;ncgen -b -o in.nc foo.cdl     note6    �      It is too troublesome to distribute in.cdl with references to NaNs because users always build with old netCDF versions that do not support it. So just comment out nan's for now.     _FillValue                              �?          FHDB �          ;J
       tm_365_�     !      tm_366�     "      tm_grg�     #      tm_jln��     $      tm_std�     %      tpt�     &      tpt_dblH�     '      tpt_fltX�     (      twod�     )      two_dmn_rec_varp�     *      two_dmn_rec_var_sng��     +      two_dmn_var��     ,      tx��     -      txyz��     .      tyت     /      tz�     1      upk��     2      upk_arr�     3      v��     4      val_eminusten��     5      val_half�     6      val_half_half��     7      val_max_max_sht	�     8      val_one_int�     9      val_one_mss!�     :      val_one_mss_int:�     ;      val_one_one_intF�     <      
var_1D_rctR�     =      
var_1D_rrg^�     >      
var_2D_rctj�     ?      
var_2D_rrgv�     @      var_msk��     A      var_nm-dash��     B      vld_rng��     C      weight��     D      wgt_one��     E      wnd_spd��     F      wvl?�     G      z��     H      zero��     I      bnd��     J      date_dmn*�     K      char_dmn_lng26n�     L      char_dmn_lng80��     M      gds_ncd��     N      vrt_nbr:�     O      char_dmn_lng04~�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          FHDB �         ���      rec_var_flt_mss_val_fltyn           rec_var_flt_mss_val_flt_all�o           #rec_var_flt_mss_val_flt_all_but_one+q           #rec_var_flt_mss_val_flt_all_but_two7t           rec_var_flt_mss_val_intxu           rec_var_flt_pck�v     	      rec_var_int_mss_val_dbl�x     
      rec_var_int_mss_val_fltz           rec_var_int_mss_val_intr{           rec_var_pck_scale_factor_only�|           rlevw~           rz�           
scalar_var�           scl_dbl_pck�           	short_var��           tdƆ           th�           threeK�           three_dmn_rec_varW�           three_dmn_var}�           three_dmn_var_crdՌ           three_dmn_var_dbl0�           three_dmn_var_int��           three_dmn_var_sht�           times�           	time_bndsO�           time_lon[�           time_udunitsg�           tm_360S�                   FHDB �         z��"�       one_dmn_rec_var_flt_scl�;     �       one_dmn_rec_var_mdnX=     �       one_dmn_rec_var_mdn__FillValued>     �       one_dmn_rec_var_missing_value�?     �       one_dmn_rec_var_mss_val�@     �       one_dmn_rec_var_mss_val_arr)B     �       one_dmn_rec_var_sngG     �       one_dmn_rec_var_unsorted�H     �       #one_dmn_rec_var_unsorted__FillValue�I     �       one_dmn_varK     �       pck_3�N     �       pck_5KQ     �       pck_7�S     �       pck_arr|V     �       piAX     �       prs_sfcMY     �       rec_var_dbl\Z     �       rec_var_dbl_mss_val_dbl_pckh[     �       rec_var_dbl_mss_val_dbl_pck_lng�]     �       rec_var_dbl_mss_val_dbl_upkT`     �       rec_var_dbl_mss_val_sht_pckc     �       rec_var_dbl_mss_val_sht_pck_shtUe     �       rec_var_dbl_mss_val_sht_upkg            rec_var_dbl_pck�i           rec_var_flt�k           rec_var_flt_mss_val_dbl�l             FHDB �         �
���       long_varH     �       lsd_dbl9     �       lsmlev�     �       masku     �       md5_a�     �       md5_abc�     �       msk_prt_mss_prt�     �       mss_val     �       mss_val_all     �       mss_val_fst)     �       mss_val_sclB     �       nan_arrN     �       nan_scl�!     �       nbdate%%     �       negative_one1(     �       nm_pnd=)     �       nm_spcI*     �       
no_mss_valU+     �       non_nul_trm_char_one_dmna,     �       non_nul_trm_char_two_dmny-     �       non_rec_var_flt_pck�.     �       od`0     �       onel1     �       one_dmn_int_val_onex2     �       one_dmn_int_val_two�3     �       one_dmn_rec_var�4     �       one_dmn_rec_var__FillValue�5     �       one_dmn_rec_var_dbl7     �       one_dmn_rec_var_flt8     �       one_dmn_rec_var_flt_mss&9     �       one_dmn_rec_var_flt_mss_scl]:     �       pckL            FHDB {�           �z     CLASS          DIMENSION_SCALE      NAME          lev      _Netcdf4Dimid                     purpose    ,      Monotonically increasing coordinate pressure     units          hybrid_sigma_pressure 	    positive          down     A_var          hyam     B_var          hybm     P0_var          P0     PS_var          PS     bounds          ilev  0   REFERENCE_LIST 6     dataset        dimension                        E�              ��             !�             ��              ��              ��              _�              k�              w�              �             }�            Ռ             p�            ��            ��            ��            �            ��                                                                                                                                                                                                                  FHDB �         ��o�       hyam��      �       hybm��      �       ilev��      �       int_var��      �       lat
�      �       
lat_1D_rct��      �       
lat_1D_rrg��      �       
lat_2D_rct��      �       
lat_2D_rrg��      �       lat_T42�      �       lat_bnd!�      �       lat_cal-�      �       lat_cpy��      �       lat_gds��      �       lat_gds_ncdQ�      �       lat_grd��      �       lat_times_long�      �       lat_times_lon_nbr��      �       lat_var\�      �       lat_wgth�      �       levt�      �       lev_cpy_�      �       lev_vark�      �       lev_wgtw�      �       lon��      �       
lon_1D_rct�      �       
lon_1D_rrg�      �       
lon_2D_rct$      �       
lon_2D_rrgD     �       lon_T42b     �       lon_calv     �       lon_gds     �       lon_gds_ncd�     �       lon_grd     �       lon_wgt�	     �       lond*     �       lonf;     0      u�     FHDB �       
  /���m       Q94!�      n       Q95-�      o       Q969�      p       Q97E�      q       Q98Q�      r       Q99]�      s       QA01i�      t       QQ01u�      u       RDM��      v       area��      w       area2��      x       area_asm��      y       att_var��      z       bnd_varE�      {       byt_2D��      |       byt_3D��      }       
byt_3D_rec��      ~       byt_arr��             byte_var��      �       byte_var_negͤ        FHDB �         Oģ�W       Q72s      X       Q73%t      Y       Q741u      Z       Q75=v      [       Q76Iw      \       Q77Uz      ]       Q78a{      ^       Q79m|      _       Q80y}      `       Q81�~      a       Q82�      b       Q83��      c       Q84��      d       Q85��      e       Q86��      f       Q87͆      g       Q88ه      h       Q89�      i       Q90�      j       Q91��      k       Q92	�      l       Q93�             FHDB �         �[UA       Q50Z      B       Q51[      C       Q52)\      D       Q535_      E       Q54A`      F       Q55Ma      G       Q56Yb      H       Q57ec      I       Q58qd      J       Q59}e      K       Q60�f      L       Q61�g      M       Q62�h      N       Q63�i      O       Q64�j      P       Q65�k      Q       Q66�l      R       Q67�m      S       Q68�n      T       Q69�o      U       Q70q      V       Q71r             FHDB �         �o�+       Q28	?      ,       Q29@      -       Q30!A      .       Q31-F      /       Q329G      0       Q33EH      1       Q34QI      2       Q35]J      3       Q36iK      4       Q37uL      5       Q38�M      6       Q39�N      7       Q40�O      8       Q41�P      9       Q42�Q      :       Q43�R      ;       Q44�S      <       Q45�T      =       Q46�U      >       Q47�V      ?       Q48�W      @       Q49Y             FHDB �         �?�       Q08$             Q09%             Q1&             Q10%'             Q1001(             Q11=)             Q12I*             Q13U+             Q14a,             Q15m-             Q16y.              Q17�/      !       Q18�0      "       Q19�5      #       Q20�6      $       Q21�7      %       Q22�8      &       Q23�9      '       Q24�:      (       Q25�;      )       Q26�<      *       Q27�=             FHDB �          VҺ        AQ01�             H2O             H2OH2OT             H2O_ice�             H2O_lqd�             H2SO4C
             Lat�             LatLon�             Lon�      	       OROD      
       P0z             PS�             Q�             Q01�             Q01Q�             Q02�             Q03�             Q04�             Q05�              Q06�!             Q07�"                     Η@{  �?  �?  �?  �?  �?     �F�     �F@              �?       @      @      @      @      @      @     �f�     �V�             �V@      �?          �?  �?       @ P�GΗ@{  �?Η@{   @  @@  �@  �@  �@  �@   A  AΗ@{   A  �B  0A  @A  PA  `A  pA  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A   B  B  B  B  B  B  B  B   B  $B  (B  ,B  0B  4B  8B  <B  @B  DB  HB  LB  PB  TB  XB  \B  `B  dB  hB  lB  pB  tB  xB  |B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �BΗ@{Η@{   A   A  �A  �@  �?   @                    	
 z�z0 ͌�C���Cf��C3��C ��C�̈C�وCf�C�           	     �B  �B      $@      $@  �B  �B  �B�_�
�@T�-@ab3/home/zender/nco/data/in.cdl                                                    /data/zender/dstccm04/dstccm04_8589_01.nc                                       /data/zender/dstccm04/dstccm04_8589_02.nc                                       /data/zender/dstccm04/dstccm04_8589_03.nc                                         �B �y�  �B �y�  �B �y�  �B �y�   A  �@��A      �?   @  @@  �@  �@  �@  �@͌�C���Cf��C3��C ��C�̈C�وCf�C͌�C���Cf��C3��C ��C�̈C�وCf�C   A   AD���l1��6�����Ky��!���P��K��¼'��@&{���o�d�0�Y���N�IWC��-8�L-���!�?�´��'^ �/i�����½��o������u���H�;F��?����k���k��?�@�?�@;FA��HA�uA��A�o�A�½A�A/i�A'^ B��B?�B��!BL-B�-8BIWCB��NB0�YB��dB��oB@&{B�'�BK��B�P�B!�BKy�B�B6��Bl1�BD��Bw^�=T3=    ��<H7�>Q~?      �C  �C �;D �;D P}D
     ��  �B  ��  ��  ��  ��  �B  �B  �B  �B  ��  ��  ��          �A  �A  �B  ��  ��  ��  ��  �B  �B  �B  �B  ��  ��  ��          �A  �A  �B�z��U/�¼������5y���¾P��F��¸'��:&{���o�d�.�Y¿�N�HWC��-8�K-���!�>�³��&^ �.i�����½��o������u���H�:F��?����k���k��?�@�?�@:FA��HA�uA��A�o�A�½A�A.i�A&^ B��B>�B��!BK-B�-8BHWCB��NB.�YB��dB��oB:&{B�'�BF��B�P�B�B5y�B��B���BU/�B�z�B  ��          �B  ��  �B     �V�      >�      >�                      >@      >@     �V@   TREE  ����������������@                                      �-             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            TREE  ����������������(                       �.             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �.             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������P                                       /             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            TREE  ����������������(                       h/             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �/             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �/             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �/             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������                              0             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             TREE  ����������������                               1             
       P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      TREE  �����������������                                              �b             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           TREE  ����������������@                              ,4             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �?       @      @      @      @      @      @       @      "@      $@     �V�      >�      >�                      >@      >@     �V@  ��      �B                           �?   @  �?   @  �B  �C  zD  �B  �C  zD  �B  �C  zD   A   @  �?      �B  4C  �C      �B  4C  �C      �B  4C  �C          4C      4C      4C          �B  4C  �C      �B  4C  �C          4C      4C      4C          4@  �@  A  4A  aA  �A ��A  �A ��A  �A ��A  B @B �B �(B  4B @?B �JB �UB  aB @lB �wB `�B  �B ��B @�B ��B ��B  �B ��B `�B  �B ��B @�B ��B ��B  �B ��B `�B  �B ��B @�B ��B ��B  �B `C 0C  C �	C �C pC @C C �C �C �C P C  #C �%C �(C �+C `.C 01C  4C �6C �9C p<C @?C BC �DC �GC �JC PMC  PC �RC �UC �XC `[C 0^C  aC �cC �fC piC @lC oC �qC �tC �wC PzC  }C �C `�C ȂC 0�C ��C  �C h�C ЉC 8�C ��C �C p�C ؐC @�C ��C �C x�C ��C H�C ��C �C ��C �C P�C ��C  �C ��C �C X�C ��C (�C ��C ��C `�C ȯC 0�C ��C      �?       @      @      @      @      @      @       @      "@      $@                     �f@             �f@             �f@                             �f@             �f@             �f@          4�  4B  C  aC ��C�>��&?��&?�>             �V@     �f@     �p@      �B  4C  �C
   ��L=���=��L>   ?  �?  @@      �?          �?  �?       @aabc   ?Η@{  �?Η@{  �BΗ@{  �BΗ@{Η@{Η@{Η@{Η@{ �y�  �B �y�  �BΗ@{      �B  �?��	   ��  �?  �?  �BΗ@{  �BΗ@{ab  abcdefghijkm      �?              �?   A    �   �-DT�!	@  zD  �C  �B     @�E ЄF   A�*
   @@      �?   @  @@  �@  �@  �@  �@   A  A   A  0A  @A  PA  `A  pA  �A  �A  �A  �A  �A  �A  �A  �A      �?   @  @@  @A  PA  `A  pA  �@  �@  �@  �@  �A  �A  �A  �A   A  A   A  0A  �A  �A  �A  �A    ػ*A    �*A    �*A     �M@     �M@     �M@     �M@     �M@     �M@   @  �?  �@  A  XA  �A  �A      @    ����              �?    ���@��.   ?   ?   ?hBhB     �?Η@{   ����            �?          �?  �?       @      �?          �?  �?       @      �?          �?  �?       @      �?          �?  �?       @      �?          �?  �?       @  �?   A   A  �?  �?TREE  ����������������P                       �f             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �f             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       g             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       -g             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       Ug             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       }g             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �g             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �g             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �g             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       h             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       Eh             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       mh             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �h             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �h             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������
                       �h             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �h             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       i             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������@                                      ?i             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            TREE  ����������������P                       j             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������                       �j             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �j             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������P                       k             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������                       [k             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������                       ok             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������P                       �k             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������                       �k             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �k             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       l             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       7l             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       _l             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �l             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �l             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �l             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������                       �l             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       m             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       ;m             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       cm             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������                       �m             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                               �m             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             TREE  ����������������@                                      �m             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            TREE  ����������������@                                      o             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            TREE  �����������������                                      Gp             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            TREE  ����������������@                                      �r             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            TREE  �����������������                                       t             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            TREE  ����������������P                       �t             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������P                               �t             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             TREE  �����������������                               Gu             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             TREE  ����������������(                       �u             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������P                       v             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       _v             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������x                               �v             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             TREE  ����������������                               �v             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             TREE  �����������������                               w             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             TREE  �����������������                                              �w             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           TREE  ����������������P                               }{             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             TREE  ����������������x                               �{             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             TREE  ����������������(                       E|             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       m|             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������(                       �|             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              TREE  ����������������@                                      �|             
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �75�7�5 ЄF @�E        ���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G���G   	   $   T   ~   ~   T   $   	         A��!A33#A��$A�j&A (A��)A33+A��,A
�/A	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOP  �?   @  @@  �@  �@  �@  �@   A  A   A  0A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A   B  B  B  B  B  B  B  B   B��	 ��	 ��	 ��	 ��	 -�	 .�	 /�	 0�	 1�	 2010-11-01T00:00:00.0000002010-11-01T01:00:00.0000002010-11-01T02:00:00.0000002010-11-01T03:00:00.0000002010-11-01T04:00:00.0000002010-11-01T05:00:00.0000002010-11-01T06:00:00.0000002010-11-01T07:00:00.0000002010-11-01T08:00:00.0000002010-11-01T09:00:00.000000/data/zender/dstccm04/dstccm04_8589_01.nc                                       /data/zender/dstccm04/dstccm04_8589_02.nc                                       /data/zender/dstccm04/dstccm04_8589_03.nc                                       /data/zender/dstccm04/dstccm04_8589_04.nc                                       /data/zender/dstccm04/dstccm04_8589_05.nc                                       /data/zender/dstccm04/dstccm04_8589_06.nc                                       /data/zender/dstccm04/dstccm04_8589_07.nc                                       /data/zender/dstccm04/dstccm04_8589_08.nc                                       /data/zender/dstccm04/dstccm04_8589_09.nc                                       /data/zender/dstccm04/dstccm04_8589_10.nc                                       ͌�C���Cf��C3��C ��C�̈C�وCf�C��C��Cf&�C33�C @�C�L�C�Y�Cff�C͌�C���Cf��C3��C ��C @�C�ىCf�C��C��Cf&�C33�C @�C @�C�Y�Cff�C͌�C���Cf��C3��C ��C ��C�يCf�C��C��Cf&�C33�C @�C�L�C�Y�Cff�C͌�C���Cf��C3��C ��C3�C�ًCf�C��C��Cf&�C33�C @�C3s�C�Y�Cff�C͌�C���Cf��C3��C ��C3�C�ٌCf�C��C��Cf&�C33�C @�C3s�C�Y�Cff�C    BTLF      :      �F� �    6     ��C �    5     �3
f A   +     e>� �   t     �j�� *   W     �7� �    5     �z� �   L     c��� P    :     �{L���                                                                                                                                                                                                                                                                                                                                                             BTLF 	     :       P    :      �    5      �    5      �    6      *   W      �   t      �   L      A   +     ����                                                                                                                                                                                                                                                                                                                                                                                                 BTLF      3      �F� �    6     ��C �    5     �3
f    +     e>� b   D     �j�� #   ?     �7� �    5     �z� �   \     c��� I    :     �{L���m                                                                                                                                                                                                                                                                                                                                                             BTLF 	     3       I    :      �    5      �    5      �    6      #   ?      b   D      �   \         +     �|�[                                                                                                                                                                                                                                                                                                                                                                                                 OCHK   �     
      +        _Netcdf4Dimid                �vƍOCHK   H�     
      +        _Netcdf4Dimid                r���OCHK   x�     
         +        _Netcdf4Dimid                5�nOCHK   ��            +        _Netcdf4Dimid             
   A�j:OCHK   <�     �       +        _Netcdf4Dimid                3YĂOCHK   ��     
   P      +        _Netcdf4Dimid                ��OCHK   ,�            +        _Netcdf4Dimid                f���OCHK   <�            +        _Netcdf4Dimid                ���OCHK                +        _Netcdf4Dimid                �W�hOCHK   x�             +        _Netcdf4Dimid                ��OCHK   ��             +        _Netcdf4Dimid                5�%OCHK   ��            +        _Netcdf4Dimid                M�w�OCHK   ��            +        _Netcdf4Dimid                ���yOCHK+        _Netcdf4Dimid                ��~OCHK+        _Netcdf4Dimid                ��~OCHK   ��             +        _Netcdf4Dimid                ��OCHK   �             +        _Netcdf4Dimid                ��6OCHK   <�             +        _Netcdf4Dimid                L}!�OCHK   \�             +        _Netcdf4Dimid                ���OCHK+        _Netcdf4Dimid                q���OCHK+        _Netcdf4Dimid                I��FOCHK   ��     @       +        _Netcdf4Dimid                �cU�OCHK   �     @       +        _Netcdf4Dimid                i�=OCHK+        _Netcdf4Dimid                I��FOCHK+        _Netcdf4Dimid                I��FOCHK+        _Netcdf4Dimid                2M< OCHK   L            +        _Netcdf4Dimid                �;�OCHK   X            +        _Netcdf4Dimid                s�IOCHK   t             +        _Netcdf4Dimid                G@m�OCHK   �             +        _Netcdf4Dimid                ��OCHK   �             +        _Netcdf4Dimid                ʯNLOCHK   �             +        _Netcdf4Dimid                d@�OCHK   D     @       +        _Netcdf4Dimid                ��s$OCHK   �     @       +        _Netcdf4Dimid                |�XGOCHK   �            +        _Netcdf4Dimid                ��9�OCHK   �             +        _Netcdf4Dimid                Ƈd�OCHK               +        _Netcdf4Dimid                �>vOCHK   h     
      +        _Netcdf4Dimid                �� wOCHK   4             +        _Netcdf4Dimid                �j��OCHK   U            +        _Netcdf4Dimid                �WNOCHK   X            +        _Netcdf4Dimid                <k��OCHK   h            +        _Netcdf4Dimid                ؊�OCHK   x            +        _Netcdf4Dimid                �-�OCHK   �            +        _Netcdf4Dimid                v)g�OCHK   �            +        _Netcdf4Dimid                ��OCHK   �            +        _Netcdf4Dimid                z�ٕOCHK   �            +        _Netcdf4Dimid                9�IOCHK   �'     
      +        _Netcdf4Dimid                ��OCHK   (0     
      +        _Netcdf4Dimid                �}eOCHK   X8     
      +        _Netcdf4Dimid                P�wgOCHK   �@     
      +        _Netcdf4Dimid                >��OCHK   �H     
      +        _Netcdf4Dimid                xG}�OCHK   �P     
      +        _Netcdf4Dimid                KDzbOCHK+        _Netcdf4Dimid                ��	OCHK   Ha     
      +        _Netcdf4Dimid                ��ϑOCHK   xi     
      +        _Netcdf4Dimid                Tl9�OCHK   �q     
      +        _Netcdf4Dimid                ]|K�OCHK   �y     
      +        _Netcdf4Dimid                ��DsOCHK   �     
      +        _Netcdf4Dimid                �P�OOCHK+        _Netcdf4Dimid                ��	OCHK   h�     
      +        _Netcdf4Dimid                ;�rOCHK+        _Netcdf4Dimid                ���kOCHK               +        _Netcdf4Dimid                �rY@OCHK                +        _Netcdf4Dimid                ﳚ#OCHK+        _Netcdf4Dimid                ��	OCHK   �     
      +        _Netcdf4Dimid                <�kOCHK   8�     
      +        _Netcdf4Dimid                ���OCHK   h�     
      +        _Netcdf4Dimid                �� �OCHK   ��     
      +        _Netcdf4Dimid                ����OCHK   ��     
      +        _Netcdf4Dimid                K�BWOCHK   ��     
      +        _Netcdf4Dimid                W�}�OCHK   (�     
      +        _Netcdf4Dimid                ^j$OCHK+        _Netcdf4Dimid                ��	OCHK   ��     
      +        _Netcdf4Dimid                nڼ`OCHK+        _Netcdf4Dimid                ��$OCHK   �      
      +        _Netcdf4Dimid                =�cMOCHK   	     
      +        _Netcdf4Dimid                o�-OCHK   H     
      +        _Netcdf4Dimid                .��	OCHK   x     
      +        _Netcdf4Dimid                i��OCHK   �!     
      +        _Netcdf4Dimid                ���>OCHK   �)     
      +        _Netcdf4Dimid                ���OCHK   2     
      +        _Netcdf4Dimid                B�	AOCHK   8:     
      +        _Netcdf4Dimid                �8$OCHK   hB     
      +        _Netcdf4Dimid                �c(�OCHK                +        _Netcdf4Dimid                ��\OCHK                +        _Netcdf4Dimid                ?q��OCHK   �T     
            +        _Netcdf4Dimid                Q��OCHK                +        _Netcdf4Dimid                ﳚ#OCHK   8     `       +        _Netcdf4Dimid                �K��OCHK   �     `       +        _Netcdf4Dimid                �l�lOCHK    ?      @ 4 4�  +        _Netcdf4Dimid                ]ʰNOCHK   �y     
            +        _Netcdf4Dimid                F��OCHK   Ѕ     
            +        _Netcdf4Dimid                9���OCHK                +        _Netcdf4Dimid                ?q��OCHK                +        _Netcdf4Dimid                ?q��OCHK   ��     
      +        _Netcdf4Dimid                �.ѿOCHK   �     
      +        _Netcdf4Dimid                ��OCHK   �     
      +        _Netcdf4Dimid                >%��OCHK                +        _Netcdf4Dimid                ﳚ#OCHK+        _Netcdf4Dimid                ��	OCHK   D            +        _Netcdf4Dimid                �h�OCHK                +        _Netcdf4Dimid                ?q��OCHK                +        _Netcdf4Dimid                ?q��OCHK                +        _Netcdf4Dimid                ?q��OCHK                +        _Netcdf4Dimid                ?q��OCHK   �     
      +        _Netcdf4Dimid                �F�
OCHK   d             +        _Netcdf4Dimid                ��e�OCHK   �     
      +        _Netcdf4Dimid                ���&OCHK   �            +        _Netcdf4Dimid                ��xOCHK   �            +        _Netcdf4Dimid                ׂIOCHK   �            +        _Netcdf4Dimid                ��?OCHK   �            +        _Netcdf4Dimid                W�ތOCHK   �            +        _Netcdf4Dimid                ��wOCHK   �             +        _Netcdf4Dimid                �1OCHK   �             +        _Netcdf4Dimid                ��OCHK   �             +        _Netcdf4Dimid                7�OCHK                +        _Netcdf4Dimid                KeEOCHK   4             +        _Netcdf4Dimid                �0pDOCHK   X            +        _Netcdf4Dimid                $���OCHK                +        _Netcdf4Dimid                �l�OCHK   x-            +        _Netcdf4Dimid                �pC�  �?   @  @@  �@  �@  �@  �@   A  A   A  0A  @A  PA  `A  pA  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A   B  B  B  B  B  B  B  B   B  $B  (B  ,B  0B  4B  8B  <B  @B  DB  HB  LB  PB  TB  XB  \B  `B  dB  hB  lB  pB  tB  xB  |B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B   C  C  C  C  C  C  C  C  C  	C  
C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C   C  !C  "C  #C  $C  %C  &C  'C  (C  )C  *C  +C  ,C  -C  .C  /C  0C  1C  2C  3C  4C  5C  6C  7C  8C  9C  :C  ;C  <C  =C  >C  ?C  @C  AC  BC  CC  DC  EC  FC  GC  HC  IC  JC  KC  LC  MC  NC  OC  PC  QC  RC  SC  TC  UC  VC  WC  XC  YC  ZC  [C  \C  ]C  ^C  _C  `C  aC  bC  cC  dC  eC  fC  gC  hC  iC  jC  kC  lC  mC  nC  oC  pC        �������?���Q��?�rh��|�?�St$��?|�Pk��?��~�Ϛ�?r���ۚ�?�ȑݚ�?_c97ݚ�?                      "   $   &                           	   
     �?   @  @@  �@  �@  �@  �@   A  AΗ@{  �?   @  @@  �@  �@  �@  �@   A  A   A  �?   @  @@  �@  �@  �@  �@   A  A   AΗ@{   @  @@  �@  �@  �@  �@   A  AΗ@{Η@{   @  @@  �@  �@  �@  �@   A  AΗ@{  �?   @  @@  �@  �@  �@  �@   A  A   A                  
   
   
   
      ���      ������
   
   
   ���  �?   @  @@  �@  �@  �@  �@   A  AΗ@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{  �?   @  @@  �@  �@  �@  �@   A  A   AHello Worl
                  	            Η@{  �@  �@   @   A  �?  A  �@  @@  �@  �?   @  @@  �@  �@  �@  �@   A  A   A  0A  @A  PA  `A  pA  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A   B  B  B  B  B  B  B  B   B  $B  (B  ,B  0B  4B  8B  <B  @B  DB  HB  LB  PB  TB  XB  \B  `B  dB  hB  lB  pB  tB  xB  |B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B      �?       @      @      @      @      @      @       @      "@      $@��UU�*  Vի��������  UU  �*      V����������������     8��       @      @      @      @      @      @       @     8��     8����UU�*  Vի������UU�*  Vի����     8��       @      @      @      @      @      @       @     8��     8��        	 
   �?   @  @@  �@  �@  �@  �@   A  A   AΗ@{   @  @@  �@  �@  �@  �@   AΗ@{Η@{Η@{   @  @@  �@  �@  �@  �@   AΗ@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{  �@Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{Η@{  �@Η@{Η@{Η@{Η@{   A �y�   @  @@  �@  �@  �@  �@   A �y� �y�        	 
 ���                     ���������                     ���������                     ������        	 
   �?   @  @@  �@  �@  �@  �@   A  A   A                        	   
                                             ��������������������������������!   "   #   $   %   &   '   (   )   *   +   ,   -   .   /   0   1   2   3   4   5   6   7   8   ����:   ;   <   =   >   ?   @   A   B   C   D   E   F   G   H   ����J   K   L   M   N   O   ����  �?   @  @@  �@  �@  �@  �@   A  A   A  0A  @A  PA  `A  pA  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A   B  B  B  B  B  B  B  B   B  $B  (B  ,B  0B  4B  8B  <B  @B  DB  HB  LB  PB  TB  XB  \B  `B  dB  hB  lB  pB  tB  xB  |B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B      �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@     �X�     �X�     �X�     �X�     �X�     �X�     �X�     �X�     �@@      A@     �A@      B@     �B@      C@     �C@      D@     �D@      E@     �E@      F@     �F@      G@     �G@      H@     �H@      I@     �I@      J@     �J@      K@     �K@      L@     �X�      M@     �M@      N@     �N@      O@     �O@      P@     @P@     �P@     �P@      Q@     @Q@     �Q@     �Q@      R@     �X�     �R@     �R@      S@     @S@     �S@     �S@     �X�                        	   
                     ��������������������������������                         !   "   #   $   %   &   '   (   )   ����+   ,   -   .   /   0   1   2   3   4   5   6   7   8   ����:   ;   <   ����>   ?   @   A   ����C   D   E   F   G   H   ����J   K   ����M   N   O   P           ��
                        ��" # ��% & ' ( ) * + , ��. / 0 1 2 3 4 5 6 7 8 9 : ; ��= > ? @ A B C D E F G H ����������������      �?       @      @      @      @      @      @       @      "@      $@   ?  �?  �?   @   @  `@  `@  �@  �@  �@  �@  �@  �@  �@  �@  A  A  A  A  (A      �B  4C  �C      �B  4C  �C      �B  4C  �C      �B  4C  �C      �B  4C  �C      �B  4C  �C      �B  4C  �C      �B  4C  �C      �B  4C  �C      �B  4C  �C͌�C���Cf��C3��C ��C�̈C�وCf�C3�C  �C�����q@33333q@�����q@fffffq@     q@�����q@33333q@�����q@fffffq@      q@͌�C���Cf��C3��C ��C�̈C�وCf�C3�C  �C  �?   @  @@  �?ff@  @@  �?��@  @@  �?33@  @@  �?��@  @@  �?   @  @@  �?ff&@  @@  �?��,@  @@  �?333@  @@  �?��9@  @@abcbcdcdedefefgfghghihijjklklm  �?   @  @@  �@  �@  �@  �@   A  A   A  0A  @A  PA  `A  pA  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A   B  B  B  B  B  B  B  B   B  �?   @  @@  �@  �@  �@  �@   A  A   A  0A  @A  PA  `A  pA  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A   B  B  B  B  B  B  B  B   B  $B  (B  ,B  0B  4B  8B  <B  @B  DB  HB  LB  PB  TB  XB  \B  `B  dB  hB  lB  pB  tB  xB  |B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B  �B   C  C  C  C  C  C  C  C  C  	C  
C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C   C  !C  "C  #C  $C  %C  &C  'C  (C  )C  *C  +C  ,C  -C  .C  /C  0C  1C  2C  3C  4C  5C  6C  7C  8C  9C  :C  ;C  <C  =C  >C  ?C  @C  AC  BC  CC  DC  EC  FC  GC  HC  IC  JC  KC  LC  MC  NC  OC  PC  QC  RC  SC  TC  UC  VC  WC  XC  YC  ZC  [C  \C  ]C  ^C  _C  `C  aC  bC  cC  dC  eC  fC  gC  hC  iC  jC  kC  lC  mC  nC  oC  pC  �?   @  @@  �@  �@  �@  �@   A  A   A  0A  @A  PA  `A  pA  �A  �A  �A  �A  �A  �?   @  @@  �@  �@  �@  �@   A  A   A  0A  @A  PA  `A  pA  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �A  �?      �?      �?      �?      �?          �?      �?      �?      �?      �? ��C �y�  4C  3C ��C  �C ��CΗ@{Η@� ��C �y�   ?  �?   ?  �?   ?  �?   ?   ? �y�   ?   ?   ?   ?   ?   ?   ?  �? �y�  �?   ?  �?   ?  �?   ?   ?   ? �y�   ?   ?   ?   ?  �?  �?  �?  �? �y�  �?  �?  �?   ?   ?   ?   ?   ? �y�   ?   ?   @   @   @   @   @   @ �y�   @   ?   ?   ?   ?   ?   ?   ? �y�   ?   ?   ?   ?   ?   ?   ?   ?   ?   ?   @   ?   ?   @   ?   ?FHDB ��          �2� 	    byte_att                       0 	    char_att          Sentence one.
Sentence two.
 
    short_att                       %      int_att                        I    	    long_att                        I    
    float_att                              �B     double_att  ?      @ 4 4�                     @R@     DIMENSION_LIST                              D�           D�             _Netcdf4Dimid                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   FHDB V          �b�k 	    byte_att                        ���� 	    char_att          Sentence one.
Sentence two.
 
    short_att                       %      int_att                        I    	    long_att                        I    
    float_att                              �B  �B  �B�B� �B�B�B     double_att  ?      @ 4 4�                     @R@      R@     �Q@q=
ף�Q@��Mb@Q@q=
ף Q@Y�;ۣ�P@     DIMENSION_LIST                              D�             _Netcdf4Dimid                                                                                                                                                                                                                                                                                                                                                                                                                                    