// -*-C++-*-
// Generate netCDF file with:
// ncgen -k netCDF-4 -b -o ~/nco/data/mdl.nc ~/nco/data/mdl.cdl

netcdf mdl {

 group: cesm {

  group: cesm_03 {
      :Conventions = "CF-1.5";
      :history = "yada yada yada";
      :Scenario = "Historical";
      :Model = "CESM";
      :Realization = "1";

    dimensions:
      time=4;
    variables:
      float tas1(time);
	  float tas2(time);
    data:
      tas1=272.3,272.3,272.3,272.3;
	  tas2=272.3,272.3,272.3,272.3;
 
    } // cesm_03

    
  } // cesm
  
 group: ecmwf {
    
  group: ecmwf_03 {
      :Conventions = "CF-1.5";
      :history = "yada yada yada";
      :Scenario = "Historical";
      :Model = "ECMWF";
      :Realization = "1";
      
    dimensions:
      time=4;
    variables:
      float tas1(time);
	  float tas2(time);
    data:
      tas1=273.3,273.3,273.3,273.3;
	  tas2=273.3,273.3,273.3,273.3;
      
    } // ecmwf_03
    
  group: ecmwf_04 {
      :Conventions = "CF-1.5";
      :history = "yada yada yada";
      :Scenario = "Historical";
      :Model = "ECMWF";
      :Realization = "2";
      
    dimensions:
      time=4;
    variables:
      float tas1(time);
	  float tas2(time);
    data:
      tas1=273.4,273.4,273.4,273.4;
	  tas2=273.4,273.4,273.4,273.4;
      
    } // ecmwf_04

  } // ecmwf

} // root group
