// Purpose: Generate a group file structure with common and non-common objects; pair of files are in_grp_1.cdl and in_grp_2.cdl
// Generate netCDF files with:
// ncgen -k netCDF-4 -b -o ~/nco/data/in_grp_1.nc ~/nco/data/in_grp_1.cdl
// ncgen -k netCDF-4 -b -o ~/nco/data/in_grp_2.nc ~/nco/data/in_grp_2.cdl

netcdf in_grp_2 {
  //
  //g1
  //
 group: g1 { 
  dimensions:
  lon1=4;
  variables:
    float var1(lon1);
  data:
    var1=0,1,1,0;
  } // end g1

} // end root group