// Generate netCDF file with:
// ncgen -k netCDF-4 -b -o ~/nco/data/cmip5.nc ~/nco/data/cmip5.cdl

netcdf cmip5 {
  dimensions:
  time=unlimited;
  :Collection = "CMIP5 RCP 8.5 Scenario";
 
  //
  //cesm
  //
  group: cesm { 
  variables:
  float tas(time);
  :Model = "CESM";
  data:
  tas=272,272,272,272;
  } // end cesm
  
  //
  //ecmwf
  //
  group: ecmwf { 
  variables:
  float tas(time);
  :Model = "ECMWF";
  data:
  tas=273,273,273,273;
  } // end ecmwf
  
  //
  //gfdl
  //
  group: gfdl { 
  variables:
  float tas(time);
  :Model = "GFDL";
  data:
  tas=274,274,274,274;
  } // end gfdl

} // end root group
