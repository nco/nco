// Purpose: CDL file to generate large netCDF test file for Large File Support (LFS) testing

// Usage:
// Create big.nc from big.cdl on a beefy 64-bit computer
// The file creation command will fail on all systems with insufficient RAM
// Transfer big.nc to a 32-bit system as an LFS testfile

// ncgen -b -o big.nc big.cdl
// ncgen -b -o ${DATA}/mie/big.nc ~/nco/data/big.cdl
// scp ~/nco/data/big.cdl esmf.ess.uci.edu:nco/data
// scp ~/nco/data/big.cdl sand.ess.uci.edu:nco/data

// Test 64-bit netCDF/NCO capabilities
// 32-bit machines do not work with files exceeding ~2 GB unless LFS enabled
// One billion floats are nco_typ_lng(NC_FLOAT)*10^9 = sizeof(float)*10^9 = 4*10^9 B = 4 GB

// Create 4 GB file with one variable 
// Expect this to fail on "small RAM" (~< 4 GB) machines:
// ncap -D 3 -O -s "wvl_1e9[wvl_1e9]=1.0f" ${DATA}/mie/big.nc ${DATA}/mie/big.nc
// ls -l ${DATA}/mie/big.nc

// On small-RAM machines, create 4 GB file with multiple variables instead
// This reduces peak memory usage to ~400 MB, and still tests LFS capability.
// ncap -D 3 -O -s "wvl_1e8[wvl_1e8]=1.0f" ${DATA}/mie/big.nc ${DATA}/mie/big.nc
// ncrename -D -d wvl_1e8,wvl big.nc # Rename because ncecat does not do coordinate variables
// Aggregate ten files together
// ncecat -D 3 -O -p ${DATA}/mie big.nc big.nc big.nc big.nc big.nc big.nc big.nc big.nc big.nc big.nc ${DATA}/mie/big.nc 
// ls -l ${DATA}/mie/big.nc

// Test data access:
// This is where LFS is useful
// These commands should work on 32-bit systems with LFS support even though files exceed 2 GB
// ncks -m -M -H ${DATA}/mie/big.nc | m
// ncks -H -d wvl_1e9,999999999 ${DATA}/mie/big.nc | m

// Valid CDF/netCDF files need not have any defined variable or data
// Use ncap LHS-casting to define variables with big dimensions
netcdf big {
dimensions:
// CDL file only used to supply dimension size = one billion to ncap 
// Create actual variable with ncap LHS-casting
	wvl_1e9=1000000000;
	wvl_1e8=100000000;
//variables:
//	float wvl_1e9(wvl_1e9);
//	float wvl_1e8(wvl_1e8);
//data:
//	wvl_1e9=1;
//	wvl_1e8=1;
}







