// -*-C++-*-
// Purpose: CDL file to generate netCDF4 test file for groups
// Created: 20110801 based on in.cdl

// Usage:
// NB: ncgen arguments depend on version:
// "-k netCDF-4" for netCDF >= 3.6.3, "-k hdf5" for netCDF < 3.6.3
// "-k netCDF-4 classic model" for netCDF >= 3.6.3, "-k hdf5-nc3" for netCDF < 3.6.3
// ncgen -k netCDF-4 -b -o ~/in_grp.nc ${HOME}/nco/data/in_grp.cdl
// scp ~/nco/data/in_grp.cdl givre.ess.uci.edu:nco/data
// scp ~/nco/data/in_grp.nc dust.ess.uci.edu:/var/www/html/nco
// scp dust.ess.uci.edu:/var/www/html/nco/in_grp.nc ~/nco/data

// Data constants in CDL:
// byte: 'a'
// char: "a"
// short: 1s
// int: 1 (no decimal point)
// float: 1.f (decimal point is required, f is required to distinguish from double)
// double: 1.0, 1.d, 1.0e-20 (decimal point is required, d is not required)

// NCL usage:
// id_in=addfile("/home/zender/nco/data/in_grp.nc","r")
// print(id_in)
// list_filevars(id_in)

netcdf in_grp {
dimensions:
	lat=2,lev=3,lon=4,gds_crd=8,time=unlimited;
variables:
	:Conventions = "CF-1.0";
	:history = "History global attribute.\n";
	:julian_day = 200000.04;
	:RCS_Header = "$Header: /data/zender/nco_20150216/nco/data/in_grp.cdl,v 1.15 2012-10-21 14:42:32 pvicente Exp $";

	float lat(lat);
	lat:long_name = "Latitude (typically midpoints)";
	lat:units = "degrees_north";

	float lev(lev);
	lev:purpose = "Monotonically increasing coordinate pressure";
	lev:units = "hybrid_sigma_pressure";
	lev:positive = "down";
	lev:A_var = "hyam";
	lev:B_var = "hybm";
	lev:P0_var = "P0";
	lev:PS_var = "PS";
	lev:bounds = "ilev";

	float lon(lon);
	lon:long_name = "Longitude (typically midpoints)";
	lon:units = "degrees_east";

	double time(time);

	float scl;

	int one_dmn_rec_var(time);
	one_dmn_rec_var:long_name = "one dimensional record variable";
	one_dmn_rec_var:units = "second";
        
	float area(lat);
	area:long_name = "area";
	area:units = "meter2";
	
	float gds_crd(gds_crd);
	gds_crd:long_name = "Geodesic coordinate";
	gds_crd:units = "degree";
	gds_crd:purpose = "enumerated coordinate like those that might define points in a geodesic grid";
	gds_crd:coordinates = "lat_gds lon_gds";

	float gds_var(gds_crd);
	gds_var:long_name = "Geodesic variable";
	gds_var:units = "meter";
	gds_var:purpose = "Test auxiliary coordinates like those that define geodesic grids";
	gds_var:coordinates = "lat_gds lon_gds";
	
	double lat_gds(gds_crd);
	lat_gds:long_name = "Latitude";  
	lat_gds:standard_name = "latitude";
	lat_gds:units="degree";
	lat_gds:purpose = "1-D latitude coordinate referred to by geodesic grid variables";

	double lon_gds(gds_crd);
	lon_gds:long_name = "Longitude";
	lon_gds:standard_name = "longitude";
	lon_gds:units="degree";
	lon_gds:purpose = "1-D longitude coordinate referred to by geodesic grid variables";


data:
	scl=1.0;
	lat=-90,90;
	lev=100,500,1000;
	lon=0,90,180,270;
	time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	one_dmn_rec_var=1,2,3,4,5,6,7,8,9,10;
	area=10.,10.;
	gds_crd=0,1,2,3,4,5,6,7;
	lat_gds=-90, -30,  -30,    0,   0, 30,  30,  90;
	lon_gds=  0,   0,  180,    0, 180,  0, 180,   0;

group: level_1_group_1 { 

      variables:
	float lon(lon);
	lon:long_name = "level_1_group_1 Longitude (typically midpoints)";
	lon:units = "level_1_group_1 degrees_east";
	float scl;
      data:
	lon=0,90,180,270;
	scl=1.1;

	group: level_2_group_1 { 
		variables:
			float scl;
		data:
			scl=1.1;
	} // end level_2_group_1

} // end level_1_group_1

group: level_1_group_2 { 
	variables:
		double time(time);
	float scl;
      data:
	time=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.;
	scl=1.2;
} // end level_1_group_2

group: level_1_group_3 {
	dimensions:
	  rlev=3,time2=unlimited;
	variables:
	  :level_1_group_3_global_attribute = "level_1_group_3_global_attribute";
	  float rz(rlev);
	  double time2(time2);
	  float scl;
	data:
	  time2=1.,2.,3.,4.,5.,6.,7.,8.,9.,10.,11.,12.,13.,14.,15.,16.,17.,18.,19.,20.;
	  rz=0,5000,17000;
	  scl=1.3;
} // end level_1_group_3

group: level_1_group_4 { 

	group: level_2_group_4 { 
	
		group: level_3_group_4 {  //group with 2 unlimited dimensions and coordinate variables
			dimensions:
			  time3=unlimited,time4=unlimited;
			variables:
			  double time3(time3);
			  double time4(time4);
			data:
			  time3=1.,2.,3.,4.,5.;
			  time4=1.,2.,3.,4.,5.,6.;
			} // end level_3_group_4
		} // end level_2_group_4
} // end level_1_group_4

group: level_1_group_5 { 

	group: level_2_group_5 { //group with 2 unlimited dimensions
			dimensions:
			  time5=unlimited,time6=unlimited;
	
		group: level_3_group_5 { 
			
			} // end level_3_group_5
		} // end level_2_group_5
} // end level_1_group_5

} // end root group
