// Purpose: CDL file to generate large netCDF test file

// Usage:
// ncgen -b -o tst.nc big.cdl
// ncgen -b -o ${DATA}/mie/big.nc ~/nco/data/big.cdl
// scp ~/nco/data/big.cdl esmf.ess.uci.edu:nco/data

// Test 64-bit netCDF/NCO capabilities
// 32-bit machines do not work with files exceeding ~2 GB
// One billion floats are nco_typ_lng(NC_FLOAT)*10^9 = sizeof(float)*10^9 = 4*10^9 B = 4 GB
// Create 4 GB file with one variable:
// ncap -s "wvl[wvl]=1.0f" ${DATA}/mie/big.nc ${DATA}/mie/big.nc
// ls -l ${DATA}/mie/big.nc

// Test data access:
// ncks -m -M -H ${DATA}/mie/big.nc | m
// ncks -H -d wvl,999999999 ${DATA}/mie/big.nc | m

// Valid CDF/netCDF files need not have any defined variable or data
// Use ncap LHS-casting to define variables with big dimensions
netcdf big {
dimensions:
	wvl=1000000000;
//variables:
//	float wvl(wvl);
//data:
//	wvl=1;
}







