// $Header Exp $
// ncgen -b -o tms_lng.nc tms_lng.cdl 

// Purpose: Template for long time-series
// Template yields initialize file size of ~10.5 MB with time as fixed dimension
// Processing is used to convert time fixed dimension to record dimension
// This is easier than initializing time with ~1 million floats in this file
// Final size is ~52.5MB, after other variables have been added

// Processing takes ~50s altogether:
// ncecat -O tms_lng.nc tms_lng.nc
// ncpdq -O -a time,record tms_lng.nc tms_lng.nc
// ncrename -O -v record,species_id tms_lng.nc tms_lng.nc
// ncap2 -O -s "hmdty[time]=98.3f;PCO2[time]=1.92f;PN2[time]=77.4f;w_vel[time]=14.8f;w_dir[time]=321.3f;temp[time]=23.5f;lmbda_260[time]=684.2f" tms_lng.nc tms_lng.nc

netcdf tms_lng{

dimensions:
    time=1314900; // Sample 8 fields at 1 Hz for one year = 8*86400*365 = 1314900

variables:
// Coordinates
    double time(time);

// 1-D variables of dimension time
    float PO2(time);
// Use for scalar weight
    double lat;

// Valid netCDF files need not have any defined variable or data
// Use ncap LHS-casting to define variables with big dimensions
// Define values for time later once ncap2 iteration works
data:
lat=76.917;
}
