// Purpose: Generate a group file structure with common and non-common objects; pair of files are in_grp_1.cdl and in_grp_2.cdl
// Generate netCDF files with:
// ncgen -k netCDF-4 -b -o ~/nco/data/in_grp_1.nc ~/nco/data/in_grp_1.cdl
// ncgen -k netCDF-4 -b -o ~/nco/data/in_grp_2.nc ~/nco/data/in_grp_2.cdl

netcdf in_grp_2 {

  dimensions:
  lon=4;
  
  //
  //g1
  //
 group: g1 { 
  variables:
    float var1(lon);
	float lon(lon);
  data:
    var1=2,2,2,2;
	lon=1,2,3,4;
  } // end g1
  
  //
  //g2
  //
 group: g2 { 
  variables:
    float var2(lon);
	float lon(lon);
  data:
    var2=2,2,2,2;
	lon=1,2,3,4;
  } // end g2  

} // end root group