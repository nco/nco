// -*-C++-*-
// Purpose: 
// ncpdq tests
// Generate netCDF files with:
// ncgen -k 4 -b -o ~/nco/data/in_grp_8.nc ~/nco/data/in_grp_8.cdl

netcdf in_grp_8 {
 group: g1 { 
   dimensions:
    lat=2;
    lon=3;
    time=unlimited;
    variables:
    float lat(lat);
    float lon(lon);
    double time(time);
    float snd(time,lat,lon);
    data:
    lat=1,2;
    lon=10,20,30;
    time=100,200;
    snd=1,2,3,4,5,6,7,8,9,10,11,12;
  } // end g1
  
  group: g2 { 
   dimensions:
    lat=2;
    lon=3;
    time=unlimited;
    variables:
    float lat(lat);
    float lon(lon);
    double time(time);
    float snd(time,lat,lon);
    data:
    lat=1,2;
    lon=10,20,30;
    time=100,200;
    snd=1,2,3,4,5,6,7,8,9,10,11,12;
  } // end g2
 
} // root group
