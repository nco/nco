netcdf test_utf8 {

dimensions:
  d2 = 2;
  xā = 2 ;
  㼿y = 2 ;
  Καλημέρα = 18 ;

variables:
  int 􍐪(xā, 㼿y) ;
  char Καλημέρα(Καλημέρα) ;
	Καλημέρα:units = "Καλημέρα" ;
  string s(xā);
  	string s:satt = "ΑΒΓΔΕΖΗΘΙΚΛΜΝΞΟΠΡΣΤΥΦΧΨΩ";

  string vs(d2);		

  // global attributes:
     :Gā = "ā㼿y􍐪" ;

data:
 􍐪 =
  1, 2,
  3, 4 ;

 Καλημέρα = "\316\232\316\261\316\273\316\267\316\274\341\275\263\317\201\316\261" ;

 s = "キャク", "龥";   

 vs = "Καλημέα" , "abc";

}
