// ncgen -k netCDF-4 -b -o ~/nco/data/clc.nc ~/nco/data/clc.cdl

netcdf clc {
  :Conventions = "CF-1.5";
  :history = "Tue Apr 25 12:46:10 PDT 2017: ncgen -k netCDF-4 -b -o ~/nco/data/clc.nc ~/nco/data/clc.cdl";
  :Purpose = "Demonstrate a collection of related datasets stored in hierarchical format";

  group: model { 
  :Source = "Model simulations, e.g., of temperature";
  dimensions:
  lat=2;
  lon=3;
  time=unlimited;
  variables:
  float temperature(time,lat,lon);
  double time(time); // Variable attributes omitted for clarity
  double lat(lat);
  double lon(lon);
  data:
  lat=-90,90.;
  lon=0.,120.,240.;
  temperature=273.,273.,273.,273.,273.,273.;
  time=1.;
  } // end model
  
  group: measurements_remote_sensing { 
  :Source = "Satellite measurements of same region as modelled, and on a different spatio-temporal grid";
  dimensions:
  lat=3;
  lon=4;
  time=unlimited;
  variables:
  float temperature(time,lat,lon);
  double time(time); // Variable attributes omitted for clarity
  double lat(lat);
  double lon(lon);
  data:
  lat=-90,0.,90.;
  lon=0.,90.,180.,270.;
  temperature=273.,273.,273.,273.,273.,273.,273.,273.,273.,273.,273.,273.;
  time=1.;
  } // end measurements_remote_sensing

  group: measurements_in_situ { 
  :Source = "In situ measurements, e.g., from an automated weather station with its own time-frequency";
  dimensions:
  time=unlimited;
  variables:
  float temperature_10m(time);
  double time(time); // Variable attributes omitted for clarity
  data:
  temperature_10m=271,272,273,274;
  time=1.,2.,3.,4.;
  } // end measurements_in_situ
  
} // end root group
