// $Header: /data/zender/nco_20150216/nco/bm/sml_stl.cdl,v 1.3 2005-06-15 22:55:51 mangalam Exp $
// when sent thru ncgen:
// ncgen -b -o smallsat.nc smallsat.cdl 

// this netCDF template should yeild a file size of ~112MB

// takes about 7.5 (real) sec on 900MHz/512MB a22p thinkpad, 
// most of it waiting for disk

// Valid CDF/netCDF files need not have any defined variable or data
// Use ncap LHS-casting to define variables with big dimensions
netcdf T85ipcc{
dimensions:
//real variables
    lat=2160; //180 degrees in 12ths of a degree from -90 to +90
    lon=4320; //360 degrees in 12ths of a degree
variables:
//indices
    double lat(lat);
    double lon(lon);

// 3 2D vars of dim 2160x4320
    float d2_00(lat,lon);
    float d2_01(lat,lon);
    float d2_02(lat,lon);

// 8 0D vars
    float weepy;

data:
lat=-89.917,-89.833,-89.750,-89.667,-89.583,-89.500,-89.417,-89.333,-89.250,-89.167,-89.083,-89.000,-88.917,-88.833,-88.750,-88.667,-88.583,-88.500,-88.417,-88.333,-88.250,-88.167,-88.083,-88.000,-87.917,-87.833,-87.750,-87.667,-87.583,-87.500,-87.417,-87.333,-87.250,-87.167,-87.083,-87.000,-86.917,-86.833,-86.750,-86.667,-86.583,-86.500,-86.417,-86.333,-86.250,-86.167,-86.083,-86.000,-85.917,-85.833,-85.750,-85.667,-85.583,-85.500,-85.417,-85.333,-85.250,-85.167,-85.083,-85.000,-84.917,-84.833,-84.750,-84.667,-84.583,-84.500,-84.417,-84.333,-84.250,-84.167,-84.083,-84.000,-83.917,-83.833,-83.750,-83.667,-83.583,-83.500,-83.417,-83.333,-83.250,-83.167,-83.083,-83.000,-82.917,-82.833,-82.750,-82.667,-82.583,-82.500,-82.417,-82.333,-82.250,-82.167,-82.083,-82.000,-81.917,-81.833,-81.750,-81.667,-81.583,-81.500,-81.417,-81.333,-81.250,-81.167,-81.083,-81.000,-80.917,-80.833,-80.750,-80.667,-80.583,-80.500,-80.417,-80.333,-80.250,-80.167,-80.083,-80.000,-79.917,-79.833,-79.750,-79.667,-79.583,-79.500,-79.417,-79.333,-79.250,-79.167,-79.083,-79.000,-78.917,-78.833,-78.750,-78.667,-78.583,-78.500,-78.417,-78.333,-78.250,-78.167,-78.083,-78.000,-77.917,-77.833,-77.750,-77.667,-77.583,-77.500,-77.417,-77.333,-77.250,-77.167,-77.083,-77.000,-76.917,-76.833,-76.750,-76.667,-76.583,-76.500,-76.417,-76.333,-76.250,-76.167,-76.083,-76.000,-75.917,-75.833,-75.750,-75.667,-75.583,-75.500,-75.417,-75.333,-75.250,-75.167,-75.083,-75.000,-74.917,-74.833,-74.750,-74.667,-74.583,-74.500,-74.417,-74.333,-74.250,-74.167,-74.083,-74.000,-73.917,-73.833,-73.750,-73.667,-73.583,-73.500,-73.417,-73.333,-73.250,-73.167,-73.083,-73.000,-72.917,-72.833,-72.750,-72.667,-72.583,-72.500,-72.417,-72.333,-72.250,-72.167,-72.083,-72.000,-71.917,-71.833,-71.750,-71.667,-71.583,-71.500,-71.417,-71.333,-71.250,-71.167,-71.083,-71.000,-70.917,-70.833,-70.750,-70.667,-70.583,-70.500,-70.417,-70.333,-70.250,-70.167,-70.083,-70.000,-69.917,-69.833,-69.750,-69.667,-69.583,-69.500,-69.417,-69.333,-69.250,-69.167,-69.083,-69.000,-68.917,-68.833,-68.750,-68.667,-68.583,-68.500,-68.417,-68.333,-68.250,-68.167,-68.083,-68.000,-67.917,-67.833,-67.750,-67.667,-67.583,-67.500,-67.417,-67.333,-67.250,-67.167,-67.083,-67.000,-66.917,-66.833,-66.750,-66.667,-66.583,-66.500,-66.417,-66.333,-66.250,-66.167,-66.083,-66.000,-65.917,-65.833,-65.750,-65.667,-65.583,-65.500,-65.417,-65.333,-65.250,-65.167,-65.083,-65.000,-64.917,-64.833,-64.750,-64.667,-64.583,-64.500,-64.417,-64.333,-64.250,-64.167,-64.083,-64.000,-63.917,-63.833,-63.750,-63.667,-63.583,-63.500,-63.417,-63.333,-63.250,-63.167,-63.083,-63.000,-62.917,-62.833,-62.750,-62.667,-62.583,-62.500,-62.417,-62.333,-62.250,-62.167,-62.083,-62.000,-61.917,-61.833,-61.750,-61.667,-61.583,-61.500,-61.417,-61.333,-61.250,-61.167,-61.083,-61.000,-60.917,-60.833,-60.750,-60.667,-60.583,-60.500,-60.417,-60.333,-60.250,-60.167,-60.083,-60.000,-59.917,-59.833,-59.750,-59.667,-59.583,-59.500,-59.417,-59.333,-59.250,-59.167,-59.083,-59.000,-58.917,-58.833,-58.750,-58.667,-58.583,-58.500,-58.417,-58.333,-58.250,-58.167,-58.083,-58.000,-57.917,-57.833,-57.750,-57.667,-57.583,-57.500,-57.417,-57.333,-57.250,-57.167,-57.083,-57.000,-56.917,-56.833,-56.750,-56.667,-56.583,-56.500,-56.417,-56.333,-56.250,-56.167,-56.083,-56.000,-55.917,-55.833,-55.750,-55.667,-55.583,-55.500,-55.417,-55.333,-55.250,-55.167,-55.083,-55.000,-54.917,-54.833,-54.750,-54.667,-54.583,-54.500,-54.417,-54.333,-54.250,-54.167,-54.083,-54.000,-53.917,-53.833,-53.750,-53.667,-53.583,-53.500,-53.417,-53.333,-53.250,-53.167,-53.083,-53.000,-52.917,-52.833,-52.750,-52.667,-52.583,-52.500,-52.417,-52.333,-52.250,-52.167,-52.083,-52.000,-51.917,-51.833,-51.750,-51.667,-51.583,-51.500,-51.417,-51.333,-51.250,-51.167,-51.083,-51.000,-50.917,-50.833,-50.750,-50.667,-50.583,-50.500,-50.417,-50.333,-50.250,-50.167,-50.083,-50.000,-49.917,-49.833,-49.750,-49.667,-49.583,-49.500,-49.417,-49.333,-49.250,-49.167,-49.083,-49.000,-48.917,-48.833,-48.750,-48.667,-48.583,-48.500,-48.417,-48.333,-48.250,-48.167,-48.083,-48.000,-47.917,-47.833,-47.750,-47.667,-47.583,-47.500,-47.417,-47.333,-47.250,-47.167,-47.083,-47.000,-46.917,-46.833,-46.750,-46.667,-46.583,-46.500,-46.417,-46.333,-46.250,-46.167,-46.083,-46.000,-45.917,-45.833,-45.750,-45.667,-45.583,-45.500,-45.417,-45.333,-45.250,-45.167,-45.083,-45.000,-44.917,-44.833,-44.750,-44.667,-44.583,-44.500,-44.417,-44.333,-44.250,-44.167,-44.083,-44.000,-43.917,-43.833,-43.750,-43.667,-43.583,-43.500,-43.417,-43.333,-43.250,-43.167,-43.083,-43.000,-42.917,-42.833,-42.750,-42.667,-42.583,-42.500,-42.417,-42.333,-42.250,-42.167,-42.083,-42.000,-41.917,-41.833,-41.750,-41.667,-41.583,-41.500,-41.417,-41.333,-41.250,-41.167,-41.083,-41.000,-40.917,-40.833,-40.750,-40.667,-40.583,-40.500,-40.417,-40.333,-40.250,-40.167,-40.083,-40.000,-39.917,-39.833,-39.750,-39.667,-39.583,-39.500,-39.417,-39.333,-39.250,-39.167,-39.083,-39.000,-38.917,-38.833,-38.750,-38.667,-38.583,-38.500,-38.417,-38.333,-38.250,-38.167,-38.083,-38.000,-37.917,-37.833,-37.750,-37.667,-37.583,-37.500,-37.417,-37.333,-37.250,-37.167,-37.083,-37.000,-36.917,-36.833,-36.750,-36.667,-36.583,-36.500,-36.417,-36.333,-36.250,-36.167,-36.083,-36.000,-35.917,-35.833,-35.750,-35.667,-35.583,-35.500,-35.417,-35.333,-35.250,-35.167,-35.083,-35.000,-34.917,-34.833,-34.750,-34.667,-34.583,-34.500,-34.417,-34.333,-34.250,-34.167,-34.083,-34.000,-33.917,-33.833,-33.750,-33.667,-33.583,-33.500,-33.417,-33.333,-33.250,-33.167,-33.083,-33.000,-32.917,-32.833,-32.750,-32.667,-32.583,-32.500,-32.417,-32.333,-32.250,-32.167,-32.083,-32.000,-31.917,-31.833,-31.750,-31.667,-31.583,-31.500,-31.417,-31.333,-31.250,-31.167,-31.083,-31.000,-30.917,-30.833,-30.750,-30.667,-30.583,-30.500,-30.417,-30.333,-30.250,-30.167,-30.083,-30.000,-29.917,-29.833,-29.750,-29.667,-29.583,-29.500,-29.417,-29.333,-29.250,-29.167,-29.083,-29.000,-28.917,-28.833,-28.750,-28.667,-28.583,-28.500,-28.417,-28.333,-28.250,-28.167,-28.083,-28.000,-27.917,-27.833,-27.750,-27.667,-27.583,-27.500,-27.417,-27.333,-27.250,-27.167,-27.083,-27.000,-26.917,-26.833,-26.750,-26.667,-26.583,-26.500,-26.417,-26.333,-26.250,-26.167,-26.083,-26.000,-25.917,-25.833,-25.750,-25.667,-25.583,-25.500,-25.417,-25.333,-25.250,-25.167,-25.083,-25.000,-24.917,-24.833,-24.750,-24.667,-24.583,-24.500,-24.417,-24.333,-24.250,-24.167,-24.083,-24.000,-23.917,-23.833,-23.750,-23.667,-23.583,-23.500,-23.417,-23.333,-23.250,-23.167,-23.083,-23.000,-22.917,-22.833,-22.750,-22.667,-22.583,-22.500,-22.417,-22.333,-22.250,-22.167,-22.083,-22.000,-21.917,-21.833,-21.750,-21.667,-21.583,-21.500,-21.417,-21.333,-21.250,-21.167,-21.083,-21.000,-20.917,-20.833,-20.750,-20.667,-20.583,-20.500,-20.417,-20.333,-20.250,-20.167,-20.083,-20.000,-19.917,-19.833,-19.750,-19.667,-19.583,-19.500,-19.417,-19.333,-19.250,-19.167,-19.083,-19.000,-18.917,-18.833,-18.750,-18.667,-18.583,-18.500,-18.417,-18.333,-18.250,-18.167,-18.083,-18.000,-17.917,-17.833,-17.750,-17.667,-17.583,-17.500,-17.417,-17.333,-17.250,-17.167,-17.083,-17.000,-16.917,-16.833,-16.750,-16.667,-16.583,-16.500,-16.417,-16.333,-16.250,-16.167,-16.083,-16.000,-15.917,-15.833,-15.750,-15.667,-15.583,-15.500,-15.417,-15.333,-15.250,-15.167,-15.083,-15.000,-14.917,-14.833,-14.750,-14.667,-14.583,-14.500,-14.417,-14.333,-14.250,-14.167,-14.083,-14.000,-13.917,-13.833,-13.750,-13.667,-13.583,-13.500,-13.417,-13.333,-13.250,-13.167,-13.083,-13.000,-12.917,-12.833,-12.750,-12.667,-12.583,-12.500,-12.417,-12.333,-12.250,-12.167,-12.083,-12.000,-11.917,-11.833,-11.750,-11.667,-11.583,-11.500,-11.417,-11.333,-11.250,-11.167,-11.083,-11.000,-10.917,-10.833,-10.750,-10.667,-10.583,-10.500,-10.417,-10.333,-10.250,-10.167,-10.083,-10.000,-9.917,-9.833,-9.750,-9.667,-9.583,-9.500,-9.417,-9.333,-9.250,-9.167,-9.083,-9.000,-8.917,-8.833,-8.750,-8.667,-8.583,-8.500,-8.417,-8.333,-8.250,-8.167,-8.083,-8.000,-7.917,-7.833,-7.750,-7.667,-7.583,-7.500,-7.417,-7.333,-7.250,-7.167,-7.083,-7.000,-6.917,-6.833,-6.750,-6.667,-6.583,-6.500,-6.417,-6.333,-6.250,-6.167,-6.083,-6.000,-5.917,-5.833,-5.750,-5.667,-5.583,-5.500,-5.417,-5.333,-5.250,-5.167,-5.083,-5.000,-4.917,-4.833,-4.750,-4.667,-4.583,-4.500,-4.417,-4.333,-4.250,-4.167,-4.083,-4.000,-3.917,-3.833,-3.750,-3.667,-3.583,-3.500,-3.417,-3.333,-3.250,-3.167,-3.083,-3.000,-2.917,-2.833,-2.750,-2.667,-2.583,-2.500,-2.417,-2.333,-2.250,-2.167,-2.083,-2.000,-1.917,-1.833,-1.750,-1.667,-1.583,-1.500,-1.417,-1.333,-1.250,-1.167,-1.083,-1.000,-0.917,-0.833,-0.750,-0.667,-0.583,-0.500,-0.417,-0.333,-0.250,-0.167,-0.083,-0.000,0.083,0.167,0.250,0.333,0.417,0.500,0.583,0.667,0.750,0.833,0.917,1.000,1.083,1.167,1.250,1.333,1.417,1.500,1.583,1.667,1.750,1.833,1.917,2.000,2.083,2.167,2.250,2.333,2.417,2.500,2.583,2.667,2.750,2.833,2.917,3.000,3.083,3.167,3.250,3.333,3.417,3.500,3.583,3.667,3.750,3.833,3.917,4.000,4.083,4.167,4.250,4.333,4.417,4.500,4.583,4.667,4.750,4.833,4.917,5.000,5.083,5.167,5.250,5.333,5.417,5.500,5.583,5.667,5.750,5.833,5.917,6.000,6.083,6.167,6.250,6.333,6.417,6.500,6.583,6.667,6.750,6.833,6.917,7.000,7.083,7.167,7.250,7.333,7.417,7.500,7.583,7.667,7.750,7.833,7.917,8.000,8.083,8.167,8.250,8.333,8.417,8.500,8.583,8.667,8.750,8.833,8.917,9.000,9.083,9.167,9.250,9.333,9.417,9.500,9.583,9.667,9.750,9.833,9.917,10.000,10.083,10.167,10.250,10.333,10.417,10.500,10.583,10.667,10.750,10.833,10.917,11.000,11.083,11.167,11.250,11.333,11.417,11.500,11.583,11.667,11.750,11.833,11.917,12.000,12.083,12.167,12.250,12.333,12.417,12.500,12.583,12.667,12.750,12.833,12.917,13.000,13.083,13.167,13.250,13.333,13.417,13.500,13.583,13.667,13.750,13.833,13.917,14.000,14.083,14.167,14.250,14.333,14.417,14.500,14.583,14.667,14.750,14.833,14.917,15.000,15.083,15.167,15.250,15.333,15.417,15.500,15.583,15.667,15.750,15.833,15.917,16.000,16.083,16.167,16.250,16.333,16.417,16.500,16.583,16.667,16.750,16.833,16.917,17.000,17.083,17.167,17.250,17.333,17.417,17.500,17.583,17.667,17.750,17.833,17.917,18.000,18.083,18.167,18.250,18.333,18.417,18.500,18.583,18.667,18.750,18.833,18.917,19.000,19.083,19.167,19.250,19.333,19.417,19.500,19.583,19.667,19.750,19.833,19.917,20.000,20.083,20.167,20.250,20.333,20.417,20.500,20.583,20.667,20.750,20.833,20.917,21.000,21.083,21.167,21.250,21.333,21.417,21.500,21.583,21.667,21.750,21.833,21.917,22.000,22.083,22.167,22.250,22.333,22.417,22.500,22.583,22.667,22.750,22.833,22.917,23.000,23.083,23.167,23.250,23.333,23.417,23.500,23.583,23.667,23.750,23.833,23.917,24.000,24.083,24.167,24.250,24.333,24.417,24.500,24.583,24.667,24.750,24.833,24.917,25.000,25.083,25.167,25.250,25.333,25.417,25.500,25.583,25.667,25.750,25.833,25.917,26.000,26.083,26.167,26.250,26.333,26.417,26.500,26.583,26.667,26.750,26.833,26.917,27.000,27.083,27.167,27.250,27.333,27.417,27.500,27.583,27.667,27.750,27.833,27.917,28.000,28.083,28.167,28.250,28.333,28.417,28.500,28.583,28.667,28.750,28.833,28.917,29.000,29.083,29.167,29.250,29.333,29.417,29.500,29.583,29.667,29.750,29.833,29.917,30.000,30.083,30.167,30.250,30.333,30.417,30.500,30.583,30.667,30.750,30.833,30.917,31.000,31.083,31.167,31.250,31.333,31.417,31.500,31.583,31.667,31.750,31.833,31.917,32.000,32.083,32.167,32.250,32.333,32.417,32.500,32.583,32.667,32.750,32.833,32.917,33.000,33.083,33.167,33.250,33.333,33.417,33.500,33.583,33.667,33.750,33.833,33.917,34.000,34.083,34.167,34.250,34.333,34.417,34.500,34.583,34.667,34.750,34.833,34.917,35.000,35.083,35.167,35.250,35.333,35.417,35.500,35.583,35.667,35.750,35.833,35.917,36.000,36.083,36.167,36.250,36.333,36.417,36.500,36.583,36.667,36.750,36.833,36.917,37.000,37.083,37.167,37.250,37.333,37.417,37.500,37.583,37.667,37.750,37.833,37.917,38.000,38.083,38.167,38.250,38.333,38.417,38.500,38.583,38.667,38.750,38.833,38.917,39.000,39.083,39.167,39.250,39.333,39.417,39.500,39.583,39.667,39.750,39.833,39.917,40.000,40.083,40.167,40.250,40.333,40.417,40.500,40.583,40.667,40.750,40.833,40.917,41.000,41.083,41.167,41.250,41.333,41.417,41.500,41.583,41.667,41.750,41.833,41.917,42.000,42.083,42.167,42.250,42.333,42.417,42.500,42.583,42.667,42.750,42.833,42.917,43.000,43.083,43.167,43.250,43.333,43.417,43.500,43.583,43.667,43.750,43.833,43.917,44.000,44.083,44.167,44.250,44.333,44.417,44.500,44.583,44.667,44.750,44.833,44.917,45.000,45.083,45.167,45.250,45.333,45.417,45.500,45.583,45.667,45.750,45.833,45.917,46.000,46.083,46.167,46.250,46.333,46.417,46.500,46.583,46.667,46.750,46.833,46.917,47.000,47.083,47.167,47.250,47.333,47.417,47.500,47.583,47.667,47.750,47.833,47.917,48.000,48.083,48.167,48.250,48.333,48.417,48.500,48.583,48.667,48.750,48.833,48.917,49.000,49.083,49.167,49.250,49.333,49.417,49.500,49.583,49.667,49.750,49.833,49.917,50.000,50.083,50.167,50.250,50.333,50.417,50.500,50.583,50.667,50.750,50.833,50.917,51.000,51.083,51.167,51.250,51.333,51.417,51.500,51.583,51.667,51.750,51.833,51.917,52.000,52.083,52.167,52.250,52.333,52.417,52.500,52.583,52.667,52.750,52.833,52.917,53.000,53.083,53.167,53.250,53.333,53.417,53.500,53.583,53.667,53.750,53.833,53.917,54.000,54.083,54.167,54.250,54.333,54.417,54.500,54.583,54.667,54.750,54.833,54.917,55.000,55.083,55.167,55.250,55.333,55.417,55.500,55.583,55.667,55.750,55.833,55.917,56.000,56.083,56.167,56.250,56.333,56.417,56.500,56.583,56.667,56.750,56.833,56.917,57.000,57.083,57.167,57.250,57.333,57.417,57.500,57.583,57.667,57.750,57.833,57.917,58.000,58.083,58.167,58.250,58.333,58.417,58.500,58.583,58.667,58.750,58.833,58.917,59.000,59.083,59.167,59.250,59.333,59.417,59.500,59.583,59.667,59.750,59.833,59.917,60.000,60.083,60.167,60.250,60.333,60.417,60.500,60.583,60.667,60.750,60.833,60.917,61.000,61.083,61.167,61.250,61.333,61.417,61.500,61.583,61.667,61.750,61.833,61.917,62.000,62.083,62.167,62.250,62.333,62.417,62.500,62.583,62.667,62.750,62.833,62.917,63.000,63.083,63.167,63.250,63.333,63.417,63.500,63.583,63.667,63.750,63.833,63.917,64.000,64.083,64.167,64.250,64.333,64.417,64.500,64.583,64.667,64.750,64.833,64.917,65.000,65.083,65.167,65.250,65.333,65.417,65.500,65.583,65.667,65.750,65.833,65.917,66.000,66.083,66.167,66.250,66.333,66.417,66.500,66.583,66.667,66.750,66.833,66.917,67.000,67.083,67.167,67.250,67.333,67.417,67.500,67.583,67.667,67.750,67.833,67.917,68.000,68.083,68.167,68.250,68.333,68.417,68.500,68.583,68.667,68.750,68.833,68.917,69.000,69.083,69.167,69.250,69.333,69.417,69.500,69.583,69.667,69.750,69.833,69.917,70.000,70.083,70.167,70.250,70.333,70.417,70.500,70.583,70.667,70.750,70.833,70.917,71.000,71.083,71.167,71.250,71.333,71.417,71.500,71.583,71.667,71.750,71.833,71.917,72.000,72.083,72.167,72.250,72.333,72.417,72.500,72.583,72.667,72.750,72.833,72.917,73.000,73.083,73.167,73.250,73.333,73.417,73.500,73.583,73.667,73.750,73.833,73.917,74.000,74.083,74.167,74.250,74.333,74.417,74.500,74.583,74.667,74.750,74.833,74.917,75.000,75.083,75.167,75.250,75.333,75.417,75.500,75.583,75.667,75.750,75.833,75.917,76.000,76.083,76.167,76.250,76.333,76.417,76.500,76.583,76.667,76.750,76.833,76.917,77.000,77.083,77.167,77.250,77.333,77.417,77.500,77.583,77.667,77.750,77.833,77.917,78.000,78.083,78.167,78.250,78.333,78.417,78.500,78.583,78.667,78.750,78.833,78.917,79.000,79.083,79.167,79.250,79.333,79.417,79.500,79.583,79.667,79.750,79.833,79.917,80.000,80.083,80.167,80.250,80.333,80.417,80.500,80.583,80.667,80.750,80.833,80.917,81.000,81.083,81.167,81.250,81.333,81.417,81.500,81.583,81.667,81.750,81.833,81.917,82.000,82.083,82.167,82.250,82.333,82.417,82.500,82.583,82.667,82.750,82.833,82.917,83.000,83.083,83.167,83.250,83.333,83.417,83.500,83.583,83.667,83.750,83.833,83.917,84.000,84.083,84.167,84.250,84.333,84.417,84.500,84.583,84.667,84.750,84.833,84.917,85.000,85.083,85.167,85.250,85.333,85.417,85.500,85.583,85.667,85.750,85.833,85.917,86.000,86.083,86.167,86.250,86.333,86.417,86.500,86.583,86.667,86.750,86.833,86.917,87.000,87.083,87.167,87.250,87.333,87.417,87.500,87.583,87.667,87.750,87.833,87.917,88.000,88.083,88.167,88.250,88.333,88.417,88.500,88.583,88.667,88.750,88.833,88.917,89.000,89.083,89.167,89.250,89.333,89.417,89.500,89.583,89.667,89.750,89.833,89.917,90.000;
lon=0.083,0.167,0.250,0.333,0.417,0.500,0.583,0.667,0.750,0.833,0.917,1.000,1.083,1.167,1.250,1.333,1.417,1.500,1.583,1.667,1.750,1.833,1.917,2.000,2.083,2.167,2.250,2.333,2.417,2.500,2.583,2.667,2.750,2.833,2.917,3.000,3.083,3.167,3.250,3.333,3.417,3.500,3.583,3.667,3.750,3.833,3.917,4.000,4.083,4.167,4.250,4.333,4.417,4.500,4.583,4.667,4.750,4.833,4.917,5.000,5.083,5.167,5.250,5.333,5.417,5.500,5.583,5.667,5.750,5.833,5.917,6.000,6.083,6.167,6.250,6.333,6.417,6.500,6.583,6.667,6.750,6.833,6.917,7.000,7.083,7.167,7.250,7.333,7.417,7.500,7.583,7.667,7.750,7.833,7.917,8.000,8.083,8.167,8.250,8.333,8.417,8.500,8.583,8.667,8.750,8.833,8.917,9.000,9.083,9.167,9.250,9.333,9.417,9.500,9.583,9.667,9.750,9.833,9.917,10.000,10.083,10.167,10.250,10.333,10.417,10.500,10.583,10.667,10.750,10.833,10.917,11.000,11.083,11.167,11.250,11.333,11.417,11.500,11.583,11.667,11.750,11.833,11.917,12.000,12.083,12.167,12.250,12.333,12.417,12.500,12.583,12.667,12.750,12.833,12.917,13.000,13.083,13.167,13.250,13.333,13.417,13.500,13.583,13.667,13.750,13.833,13.917,14.000,14.083,14.167,14.250,14.333,14.417,14.500,14.583,14.667,14.750,14.833,14.917,15.000,15.083,15.167,15.250,15.333,15.417,15.500,15.583,15.667,15.750,15.833,15.917,16.000,16.083,16.167,16.250,16.333,16.417,16.500,16.583,16.667,16.750,16.833,16.917,17.000,17.083,17.167,17.250,17.333,17.417,17.500,17.583,17.667,17.750,17.833,17.917,18.000,18.083,18.167,18.250,18.333,18.417,18.500,18.583,18.667,18.750,18.833,18.917,19.000,19.083,19.167,19.250,19.333,19.417,19.500,19.583,19.667,19.750,19.833,19.917,20.000,20.083,20.167,20.250,20.333,20.417,20.500,20.583,20.667,20.750,20.833,20.917,21.000,21.083,21.167,21.250,21.333,21.417,21.500,21.583,21.667,21.750,21.833,21.917,22.000,22.083,22.167,22.250,22.333,22.417,22.500,22.583,22.667,22.750,22.833,22.917,23.000,23.083,23.167,23.250,23.333,23.417,23.500,23.583,23.667,23.750,23.833,23.917,24.000,24.083,24.167,24.250,24.333,24.417,24.500,24.583,24.667,24.750,24.833,24.917,25.000,25.083,25.167,25.250,25.333,25.417,25.500,25.583,25.667,25.750,25.833,25.917,26.000,26.083,26.167,26.250,26.333,26.417,26.500,26.583,26.667,26.750,26.833,26.917,27.000,27.083,27.167,27.250,27.333,27.417,27.500,27.583,27.667,27.750,27.833,27.917,28.000,28.083,28.167,28.250,28.333,28.417,28.500,28.583,28.667,28.750,28.833,28.917,29.000,29.083,29.167,29.250,29.333,29.417,29.500,29.583,29.667,29.750,29.833,29.917,30.000,30.083,30.167,30.250,30.333,30.417,30.500,30.583,30.667,30.750,30.833,30.917,31.000,31.083,31.167,31.250,31.333,31.417,31.500,31.583,31.667,31.750,31.833,31.917,32.000,32.083,32.167,32.250,32.333,32.417,32.500,32.583,32.667,32.750,32.833,32.917,33.000,33.083,33.167,33.250,33.333,33.417,33.500,33.583,33.667,33.750,33.833,33.917,34.000,34.083,34.167,34.250,34.333,34.417,34.500,34.583,34.667,34.750,34.833,34.917,35.000,35.083,35.167,35.250,35.333,35.417,35.500,35.583,35.667,35.750,35.833,35.917,36.000,36.083,36.167,36.250,36.333,36.417,36.500,36.583,36.667,36.750,36.833,36.917,37.000,37.083,37.167,37.250,37.333,37.417,37.500,37.583,37.667,37.750,37.833,37.917,38.000,38.083,38.167,38.250,38.333,38.417,38.500,38.583,38.667,38.750,38.833,38.917,39.000,39.083,39.167,39.250,39.333,39.417,39.500,39.583,39.667,39.750,39.833,39.917,40.000,40.083,40.167,40.250,40.333,40.417,40.500,40.583,40.667,40.750,40.833,40.917,41.000,41.083,41.167,41.250,41.333,41.417,41.500,41.583,41.667,41.750,41.833,41.917,42.000,42.083,42.167,42.250,42.333,42.417,42.500,42.583,42.667,42.750,42.833,42.917,43.000,43.083,43.167,43.250,43.333,43.417,43.500,43.583,43.667,43.750,43.833,43.917,44.000,44.083,44.167,44.250,44.333,44.417,44.500,44.583,44.667,44.750,44.833,44.917,45.000,45.083,45.167,45.250,45.333,45.417,45.500,45.583,45.667,45.750,45.833,45.917,46.000,46.083,46.167,46.250,46.333,46.417,46.500,46.583,46.667,46.750,46.833,46.917,47.000,47.083,47.167,47.250,47.333,47.417,47.500,47.583,47.667,47.750,47.833,47.917,48.000,48.083,48.167,48.250,48.333,48.417,48.500,48.583,48.667,48.750,48.833,48.917,49.000,49.083,49.167,49.250,49.333,49.417,49.500,49.583,49.667,49.750,49.833,49.917,50.000,50.083,50.167,50.250,50.333,50.417,50.500,50.583,50.667,50.750,50.833,50.917,51.000,51.083,51.167,51.250,51.333,51.417,51.500,51.583,51.667,51.750,51.833,51.917,52.000,52.083,52.167,52.250,52.333,52.417,52.500,52.583,52.667,52.750,52.833,52.917,53.000,53.083,53.167,53.250,53.333,53.417,53.500,53.583,53.667,53.750,53.833,53.917,54.000,54.083,54.167,54.250,54.333,54.417,54.500,54.583,54.667,54.750,54.833,54.917,55.000,55.083,55.167,55.250,55.333,55.417,55.500,55.583,55.667,55.750,55.833,55.917,56.000,56.083,56.167,56.250,56.333,56.417,56.500,56.583,56.667,56.750,56.833,56.917,57.000,57.083,57.167,57.250,57.333,57.417,57.500,57.583,57.667,57.750,57.833,57.917,58.000,58.083,58.167,58.250,58.333,58.417,58.500,58.583,58.667,58.750,58.833,58.917,59.000,59.083,59.167,59.250,59.333,59.417,59.500,59.583,59.667,59.750,59.833,59.917,60.000,60.083,60.167,60.250,60.333,60.417,60.500,60.583,60.667,60.750,60.833,60.917,61.000,61.083,61.167,61.250,61.333,61.417,61.500,61.583,61.667,61.750,61.833,61.917,62.000,62.083,62.167,62.250,62.333,62.417,62.500,62.583,62.667,62.750,62.833,62.917,63.000,63.083,63.167,63.250,63.333,63.417,63.500,63.583,63.667,63.750,63.833,63.917,64.000,64.083,64.167,64.250,64.333,64.417,64.500,64.583,64.667,64.750,64.833,64.917,65.000,65.083,65.167,65.250,65.333,65.417,65.500,65.583,65.667,65.750,65.833,65.917,66.000,66.083,66.167,66.250,66.333,66.417,66.500,66.583,66.667,66.750,66.833,66.917,67.000,67.083,67.167,67.250,67.333,67.417,67.500,67.583,67.667,67.750,67.833,67.917,68.000,68.083,68.167,68.250,68.333,68.417,68.500,68.583,68.667,68.750,68.833,68.917,69.000,69.083,69.167,69.250,69.333,69.417,69.500,69.583,69.667,69.750,69.833,69.917,70.000,70.083,70.167,70.250,70.333,70.417,70.500,70.583,70.667,70.750,70.833,70.917,71.000,71.083,71.167,71.250,71.333,71.417,71.500,71.583,71.667,71.750,71.833,71.917,72.000,72.083,72.167,72.250,72.333,72.417,72.500,72.583,72.667,72.750,72.833,72.917,73.000,73.083,73.167,73.250,73.333,73.417,73.500,73.583,73.667,73.750,73.833,73.917,74.000,74.083,74.167,74.250,74.333,74.417,74.500,74.583,74.667,74.750,74.833,74.917,75.000,75.083,75.167,75.250,75.333,75.417,75.500,75.583,75.667,75.750,75.833,75.917,76.000,76.083,76.167,76.250,76.333,76.417,76.500,76.583,76.667,76.750,76.833,76.917,77.000,77.083,77.167,77.250,77.333,77.417,77.500,77.583,77.667,77.750,77.833,77.917,78.000,78.083,78.167,78.250,78.333,78.417,78.500,78.583,78.667,78.750,78.833,78.917,79.000,79.083,79.167,79.250,79.333,79.417,79.500,79.583,79.667,79.750,79.833,79.917,80.000,80.083,80.167,80.250,80.333,80.417,80.500,80.583,80.667,80.750,80.833,80.917,81.000,81.083,81.167,81.250,81.333,81.417,81.500,81.583,81.667,81.750,81.833,81.917,82.000,82.083,82.167,82.250,82.333,82.417,82.500,82.583,82.667,82.750,82.833,82.917,83.000,83.083,83.167,83.250,83.333,83.417,83.500,83.583,83.667,83.750,83.833,83.917,84.000,84.083,84.167,84.250,84.333,84.417,84.500,84.583,84.667,84.750,84.833,84.917,85.000,85.083,85.167,85.250,85.333,85.417,85.500,85.583,85.667,85.750,85.833,85.917,86.000,86.083,86.167,86.250,86.333,86.417,86.500,86.583,86.667,86.750,86.833,86.917,87.000,87.083,87.167,87.250,87.333,87.417,87.500,87.583,87.667,87.750,87.833,87.917,88.000,88.083,88.167,88.250,88.333,88.417,88.500,88.583,88.667,88.750,88.833,88.917,89.000,89.083,89.167,89.250,89.333,89.417,89.500,89.583,89.667,89.750,89.833,89.917,90.000,90.083,90.167,90.250,90.333,90.417,90.500,90.583,90.667,90.750,90.833,90.917,91.000,91.083,91.167,91.250,91.333,91.417,91.500,91.583,91.667,91.750,91.833,91.917,92.000,92.083,92.167,92.250,92.333,92.417,92.500,92.583,92.667,92.750,92.833,92.917,93.000,93.083,93.167,93.250,93.333,93.417,93.500,93.583,93.667,93.750,93.833,93.917,94.000,94.083,94.167,94.250,94.333,94.417,94.500,94.583,94.667,94.750,94.833,94.917,95.000,95.083,95.167,95.250,95.333,95.417,95.500,95.583,95.667,95.750,95.833,95.917,96.000,96.083,96.167,96.250,96.333,96.417,96.500,96.583,96.667,96.750,96.833,96.917,97.000,97.083,97.167,97.250,97.333,97.417,97.500,97.583,97.667,97.750,97.833,97.917,98.000,98.083,98.167,98.250,98.333,98.417,98.500,98.583,98.667,98.750,98.833,98.917,99.000,99.083,99.167,99.250,99.333,99.417,99.500,99.583,99.667,99.750,99.833,99.917,100.000,100.083,100.167,100.250,100.333,100.417,100.500,100.583,100.667,100.750,100.833,100.917,101.000,101.083,101.167,101.250,101.333,101.417,101.500,101.583,101.667,101.750,101.833,101.917,102.000,102.083,102.167,102.250,102.333,102.417,102.500,102.583,102.667,102.750,102.833,102.917,103.000,103.083,103.167,103.250,103.333,103.417,103.500,103.583,103.667,103.750,103.833,103.917,104.000,104.083,104.167,104.250,104.333,104.417,104.500,104.583,104.667,104.750,104.833,104.917,105.000,105.083,105.167,105.250,105.333,105.417,105.500,105.583,105.667,105.750,105.833,105.917,106.000,106.083,106.167,106.250,106.333,106.417,106.500,106.583,106.667,106.750,106.833,106.917,107.000,107.083,107.167,107.250,107.333,107.417,107.500,107.583,107.667,107.750,107.833,107.917,108.000,108.083,108.167,108.250,108.333,108.417,108.500,108.583,108.667,108.750,108.833,108.917,109.000,109.083,109.167,109.250,109.333,109.417,109.500,109.583,109.667,109.750,109.833,109.917,110.000,110.083,110.167,110.250,110.333,110.417,110.500,110.583,110.667,110.750,110.833,110.917,111.000,111.083,111.167,111.250,111.333,111.417,111.500,111.583,111.667,111.750,111.833,111.917,112.000,112.083,112.167,112.250,112.333,112.417,112.500,112.583,112.667,112.750,112.833,112.917,113.000,113.083,113.167,113.250,113.333,113.417,113.500,113.583,113.667,113.750,113.833,113.917,114.000,114.083,114.167,114.250,114.333,114.417,114.500,114.583,114.667,114.750,114.833,114.917,115.000,115.083,115.167,115.250,115.333,115.417,115.500,115.583,115.667,115.750,115.833,115.917,116.000,116.083,116.167,116.250,116.333,116.417,116.500,116.583,116.667,116.750,116.833,116.917,117.000,117.083,117.167,117.250,117.333,117.417,117.500,117.583,117.667,117.750,117.833,117.917,118.000,118.083,118.167,118.250,118.333,118.417,118.500,118.583,118.667,118.750,118.833,118.917,119.000,119.083,119.167,119.250,119.333,119.417,119.500,119.583,119.667,119.750,119.833,119.917,120.000,120.083,120.167,120.250,120.333,120.417,120.500,120.583,120.667,120.750,120.833,120.917,121.000,121.083,121.167,121.250,121.333,121.417,121.500,121.583,121.667,121.750,121.833,121.917,122.000,122.083,122.167,122.250,122.333,122.417,122.500,122.583,122.667,122.750,122.833,122.917,123.000,123.083,123.167,123.250,123.333,123.417,123.500,123.583,123.667,123.750,123.833,123.917,124.000,124.083,124.167,124.250,124.333,124.417,124.500,124.583,124.667,124.750,124.833,124.917,125.000,125.083,125.167,125.250,125.333,125.417,125.500,125.583,125.667,125.750,125.833,125.917,126.000,126.083,126.167,126.250,126.333,126.417,126.500,126.583,126.667,126.750,126.833,126.917,127.000,127.083,127.167,127.250,127.333,127.417,127.500,127.583,127.667,127.750,127.833,127.917,128.000,128.083,128.167,128.250,128.333,128.417,128.500,128.583,128.667,128.750,128.833,128.917,129.000,129.083,129.167,129.250,129.333,129.417,129.500,129.583,129.667,129.750,129.833,129.917,130.000,130.083,130.167,130.250,130.333,130.417,130.500,130.583,130.667,130.750,130.833,130.917,131.000,131.083,131.167,131.250,131.333,131.417,131.500,131.583,131.667,131.750,131.833,131.917,132.000,132.083,132.167,132.250,132.333,132.417,132.500,132.583,132.667,132.750,132.833,132.917,133.000,133.083,133.167,133.250,133.333,133.417,133.500,133.583,133.667,133.750,133.833,133.917,134.000,134.083,134.167,134.250,134.333,134.417,134.500,134.583,134.667,134.750,134.833,134.917,135.000,135.083,135.167,135.250,135.333,135.417,135.500,135.583,135.667,135.750,135.833,135.917,136.000,136.083,136.167,136.250,136.333,136.417,136.500,136.583,136.667,136.750,136.833,136.917,137.000,137.083,137.167,137.250,137.333,137.417,137.500,137.583,137.667,137.750,137.833,137.917,138.000,138.083,138.167,138.250,138.333,138.417,138.500,138.583,138.667,138.750,138.833,138.917,139.000,139.083,139.167,139.250,139.333,139.417,139.500,139.583,139.667,139.750,139.833,139.917,140.000,140.083,140.167,140.250,140.333,140.417,140.500,140.583,140.667,140.750,140.833,140.917,141.000,141.083,141.167,141.250,141.333,141.417,141.500,141.583,141.667,141.750,141.833,141.917,142.000,142.083,142.167,142.250,142.333,142.417,142.500,142.583,142.667,142.750,142.833,142.917,143.000,143.083,143.167,143.250,143.333,143.417,143.500,143.583,143.667,143.750,143.833,143.917,144.000,144.083,144.167,144.250,144.333,144.417,144.500,144.583,144.667,144.750,144.833,144.917,145.000,145.083,145.167,145.250,145.333,145.417,145.500,145.583,145.667,145.750,145.833,145.917,146.000,146.083,146.167,146.250,146.333,146.417,146.500,146.583,146.667,146.750,146.833,146.917,147.000,147.083,147.167,147.250,147.333,147.417,147.500,147.583,147.667,147.750,147.833,147.917,148.000,148.083,148.167,148.250,148.333,148.417,148.500,148.583,148.667,148.750,148.833,148.917,149.000,149.083,149.167,149.250,149.333,149.417,149.500,149.583,149.667,149.750,149.833,149.917,150.000,150.083,150.167,150.250,150.333,150.417,150.500,150.583,150.667,150.750,150.833,150.917,151.000,151.083,151.167,151.250,151.333,151.417,151.500,151.583,151.667,151.750,151.833,151.917,152.000,152.083,152.167,152.250,152.333,152.417,152.500,152.583,152.667,152.750,152.833,152.917,153.000,153.083,153.167,153.250,153.333,153.417,153.500,153.583,153.667,153.750,153.833,153.917,154.000,154.083,154.167,154.250,154.333,154.417,154.500,154.583,154.667,154.750,154.833,154.917,155.000,155.083,155.167,155.250,155.333,155.417,155.500,155.583,155.667,155.750,155.833,155.917,156.000,156.083,156.167,156.250,156.333,156.417,156.500,156.583,156.667,156.750,156.833,156.917,157.000,157.083,157.167,157.250,157.333,157.417,157.500,157.583,157.667,157.750,157.833,157.917,158.000,158.083,158.167,158.250,158.333,158.417,158.500,158.583,158.667,158.750,158.833,158.917,159.000,159.083,159.167,159.250,159.333,159.417,159.500,159.583,159.667,159.750,159.833,159.917,160.000,160.083,160.167,160.250,160.333,160.417,160.500,160.583,160.667,160.750,160.833,160.917,161.000,161.083,161.167,161.250,161.333,161.417,161.500,161.583,161.667,161.750,161.833,161.917,162.000,162.083,162.167,162.250,162.333,162.417,162.500,162.583,162.667,162.750,162.833,162.917,163.000,163.083,163.167,163.250,163.333,163.417,163.500,163.583,163.667,163.750,163.833,163.917,164.000,164.083,164.167,164.250,164.333,164.417,164.500,164.583,164.667,164.750,164.833,164.917,165.000,165.083,165.167,165.250,165.333,165.417,165.500,165.583,165.667,165.750,165.833,165.917,166.000,166.083,166.167,166.250,166.333,166.417,166.500,166.583,166.667,166.750,166.833,166.917,167.000,167.083,167.167,167.250,167.333,167.417,167.500,167.583,167.667,167.750,167.833,167.917,168.000,168.083,168.167,168.250,168.333,168.417,168.500,168.583,168.667,168.750,168.833,168.917,169.000,169.083,169.167,169.250,169.333,169.417,169.500,169.583,169.667,169.750,169.833,169.917,170.000,170.083,170.167,170.250,170.333,170.417,170.500,170.583,170.667,170.750,170.833,170.917,171.000,171.083,171.167,171.250,171.333,171.417,171.500,171.583,171.667,171.750,171.833,171.917,172.000,172.083,172.167,172.250,172.333,172.417,172.500,172.583,172.667,172.750,172.833,172.917,173.000,173.083,173.167,173.250,173.333,173.417,173.500,173.583,173.667,173.750,173.833,173.917,174.000,174.083,174.167,174.250,174.333,174.417,174.500,174.583,174.667,174.750,174.833,174.917,175.000,175.083,175.167,175.250,175.333,175.417,175.500,175.583,175.667,175.750,175.833,175.917,176.000,176.083,176.167,176.250,176.333,176.417,176.500,176.583,176.667,176.750,176.833,176.917,177.000,177.083,177.167,177.250,177.333,177.417,177.500,177.583,177.667,177.750,177.833,177.917,178.000,178.083,178.167,178.250,178.333,178.417,178.500,178.583,178.667,178.750,178.833,178.917,179.000,179.083,179.167,179.250,179.333,179.417,179.500,179.583,179.667,179.750,179.833,179.917,180.000,180.083,180.167,180.250,180.333,180.417,180.500,180.583,180.667,180.750,180.833,180.917,181.000,181.083,181.167,181.250,181.333,181.417,181.500,181.583,181.667,181.750,181.833,181.917,182.000,182.083,182.167,182.250,182.333,182.417,182.500,182.583,182.667,182.750,182.833,182.917,183.000,183.083,183.167,183.250,183.333,183.417,183.500,183.583,183.667,183.750,183.833,183.917,184.000,184.083,184.167,184.250,184.333,184.417,184.500,184.583,184.667,184.750,184.833,184.917,185.000,185.083,185.167,185.250,185.333,185.417,185.500,185.583,185.667,185.750,185.833,185.917,186.000,186.083,186.167,186.250,186.333,186.417,186.500,186.583,186.667,186.750,186.833,186.917,187.000,187.083,187.167,187.250,187.333,187.417,187.500,187.583,187.667,187.750,187.833,187.917,188.000,188.083,188.167,188.250,188.333,188.417,188.500,188.583,188.667,188.750,188.833,188.917,189.000,189.083,189.167,189.250,189.333,189.417,189.500,189.583,189.667,189.750,189.833,189.917,190.000,190.083,190.167,190.250,190.333,190.417,190.500,190.583,190.667,190.750,190.833,190.917,191.000,191.083,191.167,191.250,191.333,191.417,191.500,191.583,191.667,191.750,191.833,191.917,192.000,192.083,192.167,192.250,192.333,192.417,192.500,192.583,192.667,192.750,192.833,192.917,193.000,193.083,193.167,193.250,193.333,193.417,193.500,193.583,193.667,193.750,193.833,193.917,194.000,194.083,194.167,194.250,194.333,194.417,194.500,194.583,194.667,194.750,194.833,194.917,195.000,195.083,195.167,195.250,195.333,195.417,195.500,195.583,195.667,195.750,195.833,195.917,196.000,196.083,196.167,196.250,196.333,196.417,196.500,196.583,196.667,196.750,196.833,196.917,197.000,197.083,197.167,197.250,197.333,197.417,197.500,197.583,197.667,197.750,197.833,197.917,198.000,198.083,198.167,198.250,198.333,198.417,198.500,198.583,198.667,198.750,198.833,198.917,199.000,199.083,199.167,199.250,199.333,199.417,199.500,199.583,199.667,199.750,199.833,199.917,200.000,200.083,200.167,200.250,200.333,200.417,200.500,200.583,200.667,200.750,200.833,200.917,201.000,201.083,201.167,201.250,201.333,201.417,201.500,201.583,201.667,201.750,201.833,201.917,202.000,202.083,202.167,202.250,202.333,202.417,202.500,202.583,202.667,202.750,202.833,202.917,203.000,203.083,203.167,203.250,203.333,203.417,203.500,203.583,203.667,203.750,203.833,203.917,204.000,204.083,204.167,204.250,204.333,204.417,204.500,204.583,204.667,204.750,204.833,204.917,205.000,205.083,205.167,205.250,205.333,205.417,205.500,205.583,205.667,205.750,205.833,205.917,206.000,206.083,206.167,206.250,206.333,206.417,206.500,206.583,206.667,206.750,206.833,206.917,207.000,207.083,207.167,207.250,207.333,207.417,207.500,207.583,207.667,207.750,207.833,207.917,208.000,208.083,208.167,208.250,208.333,208.417,208.500,208.583,208.667,208.750,208.833,208.917,209.000,209.083,209.167,209.250,209.333,209.417,209.500,209.583,209.667,209.750,209.833,209.917,210.000,210.083,210.167,210.250,210.333,210.417,210.500,210.583,210.667,210.750,210.833,210.917,211.000,211.083,211.167,211.250,211.333,211.417,211.500,211.583,211.667,211.750,211.833,211.917,212.000,212.083,212.167,212.250,212.333,212.417,212.500,212.583,212.667,212.750,212.833,212.917,213.000,213.083,213.167,213.250,213.333,213.417,213.500,213.583,213.667,213.750,213.833,213.917,214.000,214.083,214.167,214.250,214.333,214.417,214.500,214.583,214.667,214.750,214.833,214.917,215.000,215.083,215.167,215.250,215.333,215.417,215.500,215.583,215.667,215.750,215.833,215.917,216.000,216.083,216.167,216.250,216.333,216.417,216.500,216.583,216.667,216.750,216.833,216.917,217.000,217.083,217.167,217.250,217.333,217.417,217.500,217.583,217.667,217.750,217.833,217.917,218.000,218.083,218.167,218.250,218.333,218.417,218.500,218.583,218.667,218.750,218.833,218.917,219.000,219.083,219.167,219.250,219.333,219.417,219.500,219.583,219.667,219.750,219.833,219.917,220.000,220.083,220.167,220.250,220.333,220.417,220.500,220.583,220.667,220.750,220.833,220.917,221.000,221.083,221.167,221.250,221.333,221.417,221.500,221.583,221.667,221.750,221.833,221.917,222.000,222.083,222.167,222.250,222.333,222.417,222.500,222.583,222.667,222.750,222.833,222.917,223.000,223.083,223.167,223.250,223.333,223.417,223.500,223.583,223.667,223.750,223.833,223.917,224.000,224.083,224.167,224.250,224.333,224.417,224.500,224.583,224.667,224.750,224.833,224.917,225.000,225.083,225.167,225.250,225.333,225.417,225.500,225.583,225.667,225.750,225.833,225.917,226.000,226.083,226.167,226.250,226.333,226.417,226.500,226.583,226.667,226.750,226.833,226.917,227.000,227.083,227.167,227.250,227.333,227.417,227.500,227.583,227.667,227.750,227.833,227.917,228.000,228.083,228.167,228.250,228.333,228.417,228.500,228.583,228.667,228.750,228.833,228.917,229.000,229.083,229.167,229.250,229.333,229.417,229.500,229.583,229.667,229.750,229.833,229.917,230.000,230.083,230.167,230.250,230.333,230.417,230.500,230.583,230.667,230.750,230.833,230.917,231.000,231.083,231.167,231.250,231.333,231.417,231.500,231.583,231.667,231.750,231.833,231.917,232.000,232.083,232.167,232.250,232.333,232.417,232.500,232.583,232.667,232.750,232.833,232.917,233.000,233.083,233.167,233.250,233.333,233.417,233.500,233.583,233.667,233.750,233.833,233.917,234.000,234.083,234.167,234.250,234.333,234.417,234.500,234.583,234.667,234.750,234.833,234.917,235.000,235.083,235.167,235.250,235.333,235.417,235.500,235.583,235.667,235.750,235.833,235.917,236.000,236.083,236.167,236.250,236.333,236.417,236.500,236.583,236.667,236.750,236.833,236.917,237.000,237.083,237.167,237.250,237.333,237.417,237.500,237.583,237.667,237.750,237.833,237.917,238.000,238.083,238.167,238.250,238.333,238.417,238.500,238.583,238.667,238.750,238.833,238.917,239.000,239.083,239.167,239.250,239.333,239.417,239.500,239.583,239.667,239.750,239.833,239.917,240.000,240.083,240.167,240.250,240.333,240.417,240.500,240.583,240.667,240.750,240.833,240.917,241.000,241.083,241.167,241.250,241.333,241.417,241.500,241.583,241.667,241.750,241.833,241.917,242.000,242.083,242.167,242.250,242.333,242.417,242.500,242.583,242.667,242.750,242.833,242.917,243.000,243.083,243.167,243.250,243.333,243.417,243.500,243.583,243.667,243.750,243.833,243.917,244.000,244.083,244.167,244.250,244.333,244.417,244.500,244.583,244.667,244.750,244.833,244.917,245.000,245.083,245.167,245.250,245.333,245.417,245.500,245.583,245.667,245.750,245.833,245.917,246.000,246.083,246.167,246.250,246.333,246.417,246.500,246.583,246.667,246.750,246.833,246.917,247.000,247.083,247.167,247.250,247.333,247.417,247.500,247.583,247.667,247.750,247.833,247.917,248.000,248.083,248.167,248.250,248.333,248.417,248.500,248.583,248.667,248.750,248.833,248.917,249.000,249.083,249.167,249.250,249.333,249.417,249.500,249.583,249.667,249.750,249.833,249.917,250.000,250.083,250.167,250.250,250.333,250.417,250.500,250.583,250.667,250.750,250.833,250.917,251.000,251.083,251.167,251.250,251.333,251.417,251.500,251.583,251.667,251.750,251.833,251.917,252.000,252.083,252.167,252.250,252.333,252.417,252.500,252.583,252.667,252.750,252.833,252.917,253.000,253.083,253.167,253.250,253.333,253.417,253.500,253.583,253.667,253.750,253.833,253.917,254.000,254.083,254.167,254.250,254.333,254.417,254.500,254.583,254.667,254.750,254.833,254.917,255.000,255.083,255.167,255.250,255.333,255.417,255.500,255.583,255.667,255.750,255.833,255.917,256.000,256.083,256.167,256.250,256.333,256.417,256.500,256.583,256.667,256.750,256.833,256.917,257.000,257.083,257.167,257.250,257.333,257.417,257.500,257.583,257.667,257.750,257.833,257.917,258.000,258.083,258.167,258.250,258.333,258.417,258.500,258.583,258.667,258.750,258.833,258.917,259.000,259.083,259.167,259.250,259.333,259.417,259.500,259.583,259.667,259.750,259.833,259.917,260.000,260.083,260.167,260.250,260.333,260.417,260.500,260.583,260.667,260.750,260.833,260.917,261.000,261.083,261.167,261.250,261.333,261.417,261.500,261.583,261.667,261.750,261.833,261.917,262.000,262.083,262.167,262.250,262.333,262.417,262.500,262.583,262.667,262.750,262.833,262.917,263.000,263.083,263.167,263.250,263.333,263.417,263.500,263.583,263.667,263.750,263.833,263.917,264.000,264.083,264.167,264.250,264.333,264.417,264.500,264.583,264.667,264.750,264.833,264.917,265.000,265.083,265.167,265.250,265.333,265.417,265.500,265.583,265.667,265.750,265.833,265.917,266.000,266.083,266.167,266.250,266.333,266.417,266.500,266.583,266.667,266.750,266.833,266.917,267.000,267.083,267.167,267.250,267.333,267.417,267.500,267.583,267.667,267.750,267.833,267.917,268.000,268.083,268.167,268.250,268.333,268.417,268.500,268.583,268.667,268.750,268.833,268.917,269.000,269.083,269.167,269.250,269.333,269.417,269.500,269.583,269.667,269.750,269.833,269.917,270.000,270.083,270.167,270.250,270.333,270.417,270.500,270.583,270.667,270.750,270.833,270.917,271.000,271.083,271.167,271.250,271.333,271.417,271.500,271.583,271.667,271.750,271.833,271.917,272.000,272.083,272.167,272.250,272.333,272.417,272.500,272.583,272.667,272.750,272.833,272.917,273.000,273.083,273.167,273.250,273.333,273.417,273.500,273.583,273.667,273.750,273.833,273.917,274.000,274.083,274.167,274.250,274.333,274.417,274.500,274.583,274.667,274.750,274.833,274.917,275.000,275.083,275.167,275.250,275.333,275.417,275.500,275.583,275.667,275.750,275.833,275.917,276.000,276.083,276.167,276.250,276.333,276.417,276.500,276.583,276.667,276.750,276.833,276.917,277.000,277.083,277.167,277.250,277.333,277.417,277.500,277.583,277.667,277.750,277.833,277.917,278.000,278.083,278.167,278.250,278.333,278.417,278.500,278.583,278.667,278.750,278.833,278.917,279.000,279.083,279.167,279.250,279.333,279.417,279.500,279.583,279.667,279.750,279.833,279.917,280.000,280.083,280.167,280.250,280.333,280.417,280.500,280.583,280.667,280.750,280.833,280.917,281.000,281.083,281.167,281.250,281.333,281.417,281.500,281.583,281.667,281.750,281.833,281.917,282.000,282.083,282.167,282.250,282.333,282.417,282.500,282.583,282.667,282.750,282.833,282.917,283.000,283.083,283.167,283.250,283.333,283.417,283.500,283.583,283.667,283.750,283.833,283.917,284.000,284.083,284.167,284.250,284.333,284.417,284.500,284.583,284.667,284.750,284.833,284.917,285.000,285.083,285.167,285.250,285.333,285.417,285.500,285.583,285.667,285.750,285.833,285.917,286.000,286.083,286.167,286.250,286.333,286.417,286.500,286.583,286.667,286.750,286.833,286.917,287.000,287.083,287.167,287.250,287.333,287.417,287.500,287.583,287.667,287.750,287.833,287.917,288.000,288.083,288.167,288.250,288.333,288.417,288.500,288.583,288.667,288.750,288.833,288.917,289.000,289.083,289.167,289.250,289.333,289.417,289.500,289.583,289.667,289.750,289.833,289.917,290.000,290.083,290.167,290.250,290.333,290.417,290.500,290.583,290.667,290.750,290.833,290.917,291.000,291.083,291.167,291.250,291.333,291.417,291.500,291.583,291.667,291.750,291.833,291.917,292.000,292.083,292.167,292.250,292.333,292.417,292.500,292.583,292.667,292.750,292.833,292.917,293.000,293.083,293.167,293.250,293.333,293.417,293.500,293.583,293.667,293.750,293.833,293.917,294.000,294.083,294.167,294.250,294.333,294.417,294.500,294.583,294.667,294.750,294.833,294.917,295.000,295.083,295.167,295.250,295.333,295.417,295.500,295.583,295.667,295.750,295.833,295.917,296.000,296.083,296.167,296.250,296.333,296.417,296.500,296.583,296.667,296.750,296.833,296.917,297.000,297.083,297.167,297.250,297.333,297.417,297.500,297.583,297.667,297.750,297.833,297.917,298.000,298.083,298.167,298.250,298.333,298.417,298.500,298.583,298.667,298.750,298.833,298.917,299.000,299.083,299.167,299.250,299.333,299.417,299.500,299.583,299.667,299.750,299.833,299.917,300.000,300.083,300.167,300.250,300.333,300.417,300.500,300.583,300.667,300.750,300.833,300.917,301.000,301.083,301.167,301.250,301.333,301.417,301.500,301.583,301.667,301.750,301.833,301.917,302.000,302.083,302.167,302.250,302.333,302.417,302.500,302.583,302.667,302.750,302.833,302.917,303.000,303.083,303.167,303.250,303.333,303.417,303.500,303.583,303.667,303.750,303.833,303.917,304.000,304.083,304.167,304.250,304.333,304.417,304.500,304.583,304.667,304.750,304.833,304.917,305.000,305.083,305.167,305.250,305.333,305.417,305.500,305.583,305.667,305.750,305.833,305.917,306.000,306.083,306.167,306.250,306.333,306.417,306.500,306.583,306.667,306.750,306.833,306.917,307.000,307.083,307.167,307.250,307.333,307.417,307.500,307.583,307.667,307.750,307.833,307.917,308.000,308.083,308.167,308.250,308.333,308.417,308.500,308.583,308.667,308.750,308.833,308.917,309.000,309.083,309.167,309.250,309.333,309.417,309.500,309.583,309.667,309.750,309.833,309.917,310.000,310.083,310.167,310.250,310.333,310.417,310.500,310.583,310.667,310.750,310.833,310.917,311.000,311.083,311.167,311.250,311.333,311.417,311.500,311.583,311.667,311.750,311.833,311.917,312.000,312.083,312.167,312.250,312.333,312.417,312.500,312.583,312.667,312.750,312.833,312.917,313.000,313.083,313.167,313.250,313.333,313.417,313.500,313.583,313.667,313.750,313.833,313.917,314.000,314.083,314.167,314.250,314.333,314.417,314.500,314.583,314.667,314.750,314.833,314.917,315.000,315.083,315.167,315.250,315.333,315.417,315.500,315.583,315.667,315.750,315.833,315.917,316.000,316.083,316.167,316.250,316.333,316.417,316.500,316.583,316.667,316.750,316.833,316.917,317.000,317.083,317.167,317.250,317.333,317.417,317.500,317.583,317.667,317.750,317.833,317.917,318.000,318.083,318.167,318.250,318.333,318.417,318.500,318.583,318.667,318.750,318.833,318.917,319.000,319.083,319.167,319.250,319.333,319.417,319.500,319.583,319.667,319.750,319.833,319.917,320.000,320.083,320.167,320.250,320.333,320.417,320.500,320.583,320.667,320.750,320.833,320.917,321.000,321.083,321.167,321.250,321.333,321.417,321.500,321.583,321.667,321.750,321.833,321.917,322.000,322.083,322.167,322.250,322.333,322.417,322.500,322.583,322.667,322.750,322.833,322.917,323.000,323.083,323.167,323.250,323.333,323.417,323.500,323.583,323.667,323.750,323.833,323.917,324.000,324.083,324.167,324.250,324.333,324.417,324.500,324.583,324.667,324.750,324.833,324.917,325.000,325.083,325.167,325.250,325.333,325.417,325.500,325.583,325.667,325.750,325.833,325.917,326.000,326.083,326.167,326.250,326.333,326.417,326.500,326.583,326.667,326.750,326.833,326.917,327.000,327.083,327.167,327.250,327.333,327.417,327.500,327.583,327.667,327.750,327.833,327.917,328.000,328.083,328.167,328.250,328.333,328.417,328.500,328.583,328.667,328.750,328.833,328.917,329.000,329.083,329.167,329.250,329.333,329.417,329.500,329.583,329.667,329.750,329.833,329.917,330.000,330.083,330.167,330.250,330.333,330.417,330.500,330.583,330.667,330.750,330.833,330.917,331.000,331.083,331.167,331.250,331.333,331.417,331.500,331.583,331.667,331.750,331.833,331.917,332.000,332.083,332.167,332.250,332.333,332.417,332.500,332.583,332.667,332.750,332.833,332.917,333.000,333.083,333.167,333.250,333.333,333.417,333.500,333.583,333.667,333.750,333.833,333.917,334.000,334.083,334.167,334.250,334.333,334.417,334.500,334.583,334.667,334.750,334.833,334.917,335.000,335.083,335.167,335.250,335.333,335.417,335.500,335.583,335.667,335.750,335.833,335.917,336.000,336.083,336.167,336.250,336.333,336.417,336.500,336.583,336.667,336.750,336.833,336.917,337.000,337.083,337.167,337.250,337.333,337.417,337.500,337.583,337.667,337.750,337.833,337.917,338.000,338.083,338.167,338.250,338.333,338.417,338.500,338.583,338.667,338.750,338.833,338.917,339.000,339.083,339.167,339.250,339.333,339.417,339.500,339.583,339.667,339.750,339.833,339.917,340.000,340.083,340.167,340.250,340.333,340.417,340.500,340.583,340.667,340.750,340.833,340.917,341.000,341.083,341.167,341.250,341.333,341.417,341.500,341.583,341.667,341.750,341.833,341.917,342.000,342.083,342.167,342.250,342.333,342.417,342.500,342.583,342.667,342.750,342.833,342.917,343.000,343.083,343.167,343.250,343.333,343.417,343.500,343.583,343.667,343.750,343.833,343.917,344.000,344.083,344.167,344.250,344.333,344.417,344.500,344.583,344.667,344.750,344.833,344.917,345.000,345.083,345.167,345.250,345.333,345.417,345.500,345.583,345.667,345.750,345.833,345.917,346.000,346.083,346.167,346.250,346.333,346.417,346.500,346.583,346.667,346.750,346.833,346.917,347.000,347.083,347.167,347.250,347.333,347.417,347.500,347.583,347.667,347.750,347.833,347.917,348.000,348.083,348.167,348.250,348.333,348.417,348.500,348.583,348.667,348.750,348.833,348.917,349.000,349.083,349.167,349.250,349.333,349.417,349.500,349.583,349.667,349.750,349.833,349.917,350.000,350.083,350.167,350.250,350.333,350.417,350.500,350.583,350.667,350.750,350.833,350.917,351.000,351.083,351.167,351.250,351.333,351.417,351.500,351.583,351.667,351.750,351.833,351.917,352.000,352.083,352.167,352.250,352.333,352.417,352.500,352.583,352.667,352.750,352.833,352.917,353.000,353.083,353.167,353.250,353.333,353.417,353.500,353.583,353.667,353.750,353.833,353.917,354.000,354.083,354.167,354.250,354.333,354.417,354.500,354.583,354.667,354.750,354.833,354.917,355.000,355.083,355.167,355.250,355.333,355.417,355.500,355.583,355.667,355.750,355.833,355.917,356.000,356.083,356.167,356.250,356.333,356.417,356.500,356.583,356.667,356.750,356.833,356.917,357.000,357.083,357.167,357.250,357.333,357.417,357.500,357.583,357.667,357.750,357.833,357.917,358.000,358.083,358.167,358.250,358.333,358.417,358.500,358.583,358.667,358.750,358.833,358.917,359.000,359.083,359.167,359.250,359.333,359.417,359.500,359.583,359.667,359.750,359.833,359.917, 360.000;
weepy=1.23456;
}
